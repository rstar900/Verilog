// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jul 24 2022 20:50:09

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "led_blink_top" view "INTERFACE"

module led_blink_top (
    o_LED_3,
    o_LED_1,
    i_Clk,
    o_LED_4,
    o_LED_2);

    output o_LED_3;
    output o_LED_1;
    input i_Clk;
    output o_LED_4;
    output o_LED_2;

    wire N__5323;
    wire N__5322;
    wire N__5321;
    wire N__5312;
    wire N__5311;
    wire N__5310;
    wire N__5303;
    wire N__5302;
    wire N__5301;
    wire N__5294;
    wire N__5293;
    wire N__5292;
    wire N__5285;
    wire N__5284;
    wire N__5283;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5245;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5233;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5215;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5191;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5176;
    wire N__5175;
    wire N__5174;
    wire N__5171;
    wire N__5170;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5152;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5142;
    wire N__5137;
    wire N__5136;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5113;
    wire N__5110;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5098;
    wire N__5095;
    wire N__5092;
    wire N__5091;
    wire N__5090;
    wire N__5089;
    wire N__5088;
    wire N__5087;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5079;
    wire N__5078;
    wire N__5073;
    wire N__5062;
    wire N__5057;
    wire N__5054;
    wire N__5047;
    wire N__5046;
    wire N__5041;
    wire N__5040;
    wire N__5039;
    wire N__5038;
    wire N__5037;
    wire N__5036;
    wire N__5035;
    wire N__5034;
    wire N__5031;
    wire N__5022;
    wire N__5015;
    wire N__5008;
    wire N__5005;
    wire N__5002;
    wire N__4999;
    wire N__4998;
    wire N__4995;
    wire N__4994;
    wire N__4993;
    wire N__4992;
    wire N__4991;
    wire N__4990;
    wire N__4989;
    wire N__4984;
    wire N__4983;
    wire N__4982;
    wire N__4979;
    wire N__4968;
    wire N__4965;
    wire N__4958;
    wire N__4951;
    wire N__4950;
    wire N__4949;
    wire N__4948;
    wire N__4947;
    wire N__4946;
    wire N__4945;
    wire N__4944;
    wire N__4943;
    wire N__4942;
    wire N__4941;
    wire N__4940;
    wire N__4939;
    wire N__4938;
    wire N__4937;
    wire N__4936;
    wire N__4935;
    wire N__4934;
    wire N__4933;
    wire N__4932;
    wire N__4931;
    wire N__4930;
    wire N__4929;
    wire N__4928;
    wire N__4927;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4855;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4845;
    wire N__4840;
    wire N__4839;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4825;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4789;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4777;
    wire N__4774;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4762;
    wire N__4761;
    wire N__4758;
    wire N__4755;
    wire N__4750;
    wire N__4749;
    wire N__4746;
    wire N__4743;
    wire N__4740;
    wire N__4735;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4723;
    wire N__4722;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4705;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4669;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4657;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4645;
    wire N__4644;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4630;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4618;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4573;
    wire N__4570;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4560;
    wire N__4555;
    wire N__4552;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4537;
    wire N__4534;
    wire N__4531;
    wire N__4528;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4417;
    wire N__4414;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4399;
    wire N__4396;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4360;
    wire N__4357;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4342;
    wire N__4339;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4324;
    wire N__4321;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4300;
    wire N__4297;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4285;
    wire N__4282;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4270;
    wire N__4267;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4257;
    wire N__4252;
    wire N__4249;
    wire N__4248;
    wire N__4245;
    wire N__4242;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4186;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4113;
    wire N__4112;
    wire N__4107;
    wire N__4104;
    wire N__4099;
    wire N__4098;
    wire N__4097;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4085;
    wire N__4082;
    wire N__4075;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4060;
    wire N__4057;
    wire N__4054;
    wire N__4051;
    wire N__4048;
    wire N__4045;
    wire N__4042;
    wire N__4041;
    wire N__4040;
    wire N__4039;
    wire N__4038;
    wire N__4037;
    wire N__4036;
    wire N__4029;
    wire N__4028;
    wire N__4027;
    wire N__4024;
    wire N__4023;
    wire N__4016;
    wire N__4013;
    wire N__4006;
    wire N__4003;
    wire N__3994;
    wire N__3993;
    wire N__3992;
    wire N__3991;
    wire N__3990;
    wire N__3989;
    wire N__3988;
    wire N__3987;
    wire N__3986;
    wire N__3979;
    wire N__3972;
    wire N__3965;
    wire N__3958;
    wire N__3957;
    wire N__3956;
    wire N__3955;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3947;
    wire N__3946;
    wire N__3943;
    wire N__3942;
    wire N__3941;
    wire N__3938;
    wire N__3935;
    wire N__3930;
    wire N__3923;
    wire N__3916;
    wire N__3907;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3889;
    wire N__3886;
    wire N__3883;
    wire N__3880;
    wire N__3877;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3867;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3850;
    wire N__3847;
    wire N__3844;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3817;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3802;
    wire N__3801;
    wire N__3798;
    wire N__3797;
    wire N__3796;
    wire N__3795;
    wire N__3794;
    wire N__3793;
    wire N__3792;
    wire N__3791;
    wire N__3790;
    wire N__3789;
    wire N__3788;
    wire N__3787;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3767;
    wire N__3764;
    wire N__3757;
    wire N__3750;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3732;
    wire N__3731;
    wire N__3730;
    wire N__3729;
    wire N__3728;
    wire N__3727;
    wire N__3726;
    wire N__3725;
    wire N__3724;
    wire N__3723;
    wire N__3722;
    wire N__3721;
    wire N__3718;
    wire N__3705;
    wire N__3698;
    wire N__3691;
    wire N__3682;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3672;
    wire N__3671;
    wire N__3670;
    wire N__3669;
    wire N__3666;
    wire N__3665;
    wire N__3664;
    wire N__3661;
    wire N__3660;
    wire N__3657;
    wire N__3656;
    wire N__3655;
    wire N__3652;
    wire N__3651;
    wire N__3650;
    wire N__3647;
    wire N__3646;
    wire N__3643;
    wire N__3630;
    wire N__3627;
    wire N__3620;
    wire N__3615;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3595;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3583;
    wire N__3580;
    wire N__3577;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3565;
    wire N__3562;
    wire N__3561;
    wire N__3558;
    wire N__3555;
    wire N__3550;
    wire N__3547;
    wire N__3544;
    wire N__3541;
    wire N__3540;
    wire N__3537;
    wire N__3534;
    wire N__3531;
    wire N__3528;
    wire N__3523;
    wire N__3520;
    wire N__3519;
    wire N__3516;
    wire N__3513;
    wire N__3510;
    wire N__3505;
    wire N__3502;
    wire N__3499;
    wire N__3496;
    wire N__3493;
    wire N__3490;
    wire N__3489;
    wire N__3486;
    wire N__3483;
    wire N__3480;
    wire N__3475;
    wire N__3472;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3460;
    wire N__3457;
    wire N__3454;
    wire N__3453;
    wire N__3450;
    wire N__3447;
    wire N__3444;
    wire N__3439;
    wire N__3436;
    wire N__3433;
    wire N__3430;
    wire N__3427;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3417;
    wire N__3412;
    wire N__3409;
    wire N__3406;
    wire N__3403;
    wire N__3400;
    wire N__3397;
    wire N__3394;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3384;
    wire N__3379;
    wire N__3376;
    wire N__3373;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3363;
    wire N__3360;
    wire N__3357;
    wire N__3352;
    wire N__3349;
    wire N__3348;
    wire N__3345;
    wire N__3342;
    wire N__3337;
    wire N__3334;
    wire N__3333;
    wire N__3330;
    wire N__3327;
    wire N__3324;
    wire N__3319;
    wire N__3316;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3304;
    wire N__3301;
    wire N__3300;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3283;
    wire N__3280;
    wire N__3277;
    wire N__3274;
    wire N__3271;
    wire N__3270;
    wire N__3267;
    wire N__3264;
    wire N__3261;
    wire N__3256;
    wire N__3253;
    wire N__3250;
    wire N__3247;
    wire N__3244;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3231;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3210;
    wire N__3207;
    wire N__3204;
    wire N__3201;
    wire N__3198;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3184;
    wire N__3181;
    wire N__3178;
    wire N__3175;
    wire N__3172;
    wire N__3169;
    wire N__3166;
    wire N__3163;
    wire N__3160;
    wire N__3159;
    wire N__3154;
    wire N__3153;
    wire N__3150;
    wire N__3147;
    wire N__3142;
    wire N__3141;
    wire N__3138;
    wire N__3137;
    wire N__3136;
    wire N__3133;
    wire N__3126;
    wire N__3123;
    wire N__3118;
    wire N__3117;
    wire N__3114;
    wire N__3111;
    wire N__3108;
    wire N__3105;
    wire N__3100;
    wire N__3097;
    wire N__3096;
    wire N__3093;
    wire N__3090;
    wire N__3085;
    wire N__3082;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3057;
    wire N__3054;
    wire N__3051;
    wire N__3048;
    wire N__3045;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3030;
    wire N__3029;
    wire N__3028;
    wire N__3027;
    wire N__3026;
    wire N__3025;
    wire N__3024;
    wire N__3023;
    wire N__3022;
    wire N__3019;
    wire N__3010;
    wire N__2999;
    wire N__2998;
    wire N__2997;
    wire N__2996;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2977;
    wire N__2968;
    wire N__2967;
    wire N__2966;
    wire N__2965;
    wire N__2964;
    wire N__2963;
    wire N__2962;
    wire N__2961;
    wire N__2960;
    wire N__2959;
    wire N__2958;
    wire N__2957;
    wire N__2956;
    wire N__2953;
    wire N__2944;
    wire N__2935;
    wire N__2926;
    wire N__2917;
    wire N__2914;
    wire N__2913;
    wire N__2912;
    wire N__2911;
    wire N__2910;
    wire N__2909;
    wire N__2908;
    wire N__2907;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2896;
    wire N__2895;
    wire N__2892;
    wire N__2891;
    wire N__2890;
    wire N__2887;
    wire N__2884;
    wire N__2881;
    wire N__2878;
    wire N__2869;
    wire N__2860;
    wire N__2851;
    wire N__2842;
    wire N__2839;
    wire N__2836;
    wire N__2835;
    wire N__2832;
    wire N__2829;
    wire N__2824;
    wire N__2821;
    wire N__2820;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2808;
    wire N__2803;
    wire N__2800;
    wire N__2797;
    wire N__2794;
    wire N__2793;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2776;
    wire N__2773;
    wire N__2772;
    wire N__2769;
    wire N__2766;
    wire N__2763;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2728;
    wire N__2725;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2715;
    wire N__2710;
    wire N__2707;
    wire N__2704;
    wire N__2701;
    wire N__2700;
    wire N__2697;
    wire N__2694;
    wire N__2691;
    wire N__2686;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2667;
    wire N__2662;
    wire N__2659;
    wire N__2656;
    wire N__2653;
    wire N__2652;
    wire N__2649;
    wire N__2646;
    wire N__2643;
    wire N__2638;
    wire N__2635;
    wire N__2632;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2622;
    wire N__2619;
    wire N__2616;
    wire N__2613;
    wire N__2608;
    wire N__2605;
    wire N__2602;
    wire N__2599;
    wire N__2596;
    wire N__2595;
    wire N__2592;
    wire N__2589;
    wire N__2584;
    wire N__2581;
    wire N__2578;
    wire N__2575;
    wire N__2574;
    wire N__2571;
    wire N__2568;
    wire N__2563;
    wire N__2560;
    wire N__2559;
    wire N__2556;
    wire N__2553;
    wire N__2550;
    wire N__2545;
    wire N__2542;
    wire N__2541;
    wire N__2538;
    wire N__2535;
    wire N__2532;
    wire N__2527;
    wire N__2524;
    wire N__2523;
    wire N__2520;
    wire N__2517;
    wire N__2512;
    wire N__2509;
    wire N__2506;
    wire N__2503;
    wire N__2500;
    wire N__2497;
    wire N__2496;
    wire N__2493;
    wire N__2490;
    wire N__2485;
    wire N__2482;
    wire N__2479;
    wire N__2476;
    wire N__2475;
    wire N__2472;
    wire N__2469;
    wire N__2466;
    wire N__2461;
    wire N__2458;
    wire N__2455;
    wire N__2452;
    wire N__2451;
    wire N__2448;
    wire N__2445;
    wire N__2442;
    wire N__2437;
    wire N__2434;
    wire N__2431;
    wire N__2428;
    wire N__2425;
    wire N__2422;
    wire N__2421;
    wire N__2420;
    wire N__2417;
    wire N__2414;
    wire N__2411;
    wire N__2404;
    wire N__2403;
    wire N__2402;
    wire N__2401;
    wire N__2398;
    wire N__2395;
    wire N__2392;
    wire N__2389;
    wire N__2386;
    wire N__2377;
    wire N__2374;
    wire N__2373;
    wire N__2370;
    wire N__2367;
    wire N__2362;
    wire N__2359;
    wire N__2358;
    wire N__2355;
    wire N__2352;
    wire N__2347;
    wire N__2344;
    wire N__2343;
    wire N__2340;
    wire N__2337;
    wire N__2334;
    wire N__2329;
    wire N__2326;
    wire N__2325;
    wire N__2322;
    wire N__2319;
    wire N__2314;
    wire N__2311;
    wire N__2308;
    wire N__2305;
    wire N__2302;
    wire N__2299;
    wire N__2296;
    wire N__2293;
    wire N__2290;
    wire N__2287;
    wire N__2284;
    wire N__2281;
    wire N__2278;
    wire N__2275;
    wire N__2272;
    wire N__2269;
    wire N__2266;
    wire N__2265;
    wire N__2262;
    wire N__2259;
    wire VCCG0;
    wire GNDG0;
    wire o_LED_1_c;
    wire \led_blink_inst.o_LED_13_15 ;
    wire \led_blink_inst.o_LED_13_13 ;
    wire \led_blink_inst.o_LED_13_14_cascade_ ;
    wire \led_blink_inst.o_LED_13_12 ;
    wire \led_blink_inst.o_LED_13_21_cascade_ ;
    wire \led_blink_inst.o_LED_13_16_cascade_ ;
    wire \led_blink_inst.o_LED_23_16_cascade_ ;
    wire \led_blink_inst.r_Count_1Z0Z_1 ;
    wire \led_blink_inst.r_Count_1Z0Z_0 ;
    wire bfn_8_7_0_;
    wire \led_blink_inst.r_Count_1Z0Z_2 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_1 ;
    wire \led_blink_inst.r_Count_1Z0Z_3 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_2 ;
    wire \led_blink_inst.r_Count_1Z0Z_4 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_3 ;
    wire \led_blink_inst.r_Count_1Z0Z_5 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_5 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_4 ;
    wire \led_blink_inst.r_Count_1Z0Z_6 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_5 ;
    wire \led_blink_inst.r_Count_1Z0Z_7 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_6 ;
    wire \led_blink_inst.r_Count_1Z0Z_8 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_7 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_8 ;
    wire \led_blink_inst.r_Count_1Z0Z_9 ;
    wire bfn_8_8_0_;
    wire \led_blink_inst.r_Count_1Z0Z_10 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_10 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_9 ;
    wire \led_blink_inst.r_Count_1Z0Z_11 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_11 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_10 ;
    wire \led_blink_inst.r_Count_1Z0Z_12 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_12 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_11 ;
    wire \led_blink_inst.r_Count_1Z0Z_13 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_13 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_12 ;
    wire \led_blink_inst.r_Count_1Z0Z_14 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_13 ;
    wire \led_blink_inst.r_Count_1Z0Z_15 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_15 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_14 ;
    wire \led_blink_inst.r_Count_1Z0Z_16 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_15 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_16 ;
    wire \led_blink_inst.r_Count_1Z0Z_17 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_17 ;
    wire bfn_8_9_0_;
    wire \led_blink_inst.r_Count_1Z0Z_18 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_18 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_17 ;
    wire \led_blink_inst.r_Count_1Z0Z_19 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_19 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_18 ;
    wire \led_blink_inst.r_Count_1Z0Z_20 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_20 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_19 ;
    wire \led_blink_inst.r_Count_1Z0Z_21 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_21 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_20 ;
    wire \led_blink_inst.r_Count_1Z0Z_22 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_21 ;
    wire \led_blink_inst.un3_r_Count_1_1_cry_22 ;
    wire \led_blink_inst.o_LED_13_17 ;
    wire \led_blink_inst.o_LED_13_16 ;
    wire \led_blink_inst.r_Count_1_RNO_0Z0Z_23_cascade_ ;
    wire \led_blink_inst.o_LED_13_21 ;
    wire \led_blink_inst.r_Count_1Z0Z_23 ;
    wire o_LED_2_c;
    wire \led_blink_inst.o_LED_23_14 ;
    wire \led_blink_inst.o_LED_23_13 ;
    wire \led_blink_inst.o_LED_23_12_cascade_ ;
    wire \led_blink_inst.o_LED_23_15 ;
    wire \led_blink_inst.o_LED_23_21_cascade_ ;
    wire \led_blink_inst.r_Count_2Z0Z_1 ;
    wire \led_blink_inst.r_Count_2Z0Z_0 ;
    wire bfn_9_6_0_;
    wire \led_blink_inst.r_Count_2Z0Z_2 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_1 ;
    wire \led_blink_inst.r_Count_2Z0Z_3 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_2 ;
    wire \led_blink_inst.r_Count_2Z0Z_4 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_4 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_3 ;
    wire \led_blink_inst.r_Count_2Z0Z_5 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_4 ;
    wire \led_blink_inst.r_Count_2Z0Z_6 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_5 ;
    wire \led_blink_inst.r_Count_2Z0Z_7 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_6 ;
    wire \led_blink_inst.r_Count_2Z0Z_8 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_7 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_8 ;
    wire \led_blink_inst.r_Count_2Z0Z_9 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_9 ;
    wire bfn_9_7_0_;
    wire \led_blink_inst.r_Count_2Z0Z_10 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_10 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_9 ;
    wire \led_blink_inst.r_Count_2Z0Z_11 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_11 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_10 ;
    wire \led_blink_inst.r_Count_2Z0Z_12 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_12 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_11 ;
    wire \led_blink_inst.r_Count_2Z0Z_13 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_12 ;
    wire \led_blink_inst.r_Count_2Z0Z_14 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_14 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_13 ;
    wire \led_blink_inst.r_Count_2Z0Z_15 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_14 ;
    wire \led_blink_inst.r_Count_2Z0Z_16 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_16 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_15 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_16 ;
    wire \led_blink_inst.r_Count_2Z0Z_17 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_17 ;
    wire bfn_9_8_0_;
    wire \led_blink_inst.r_Count_2Z0Z_18 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_18 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_17 ;
    wire \led_blink_inst.r_Count_2Z0Z_19 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_19 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_18 ;
    wire \led_blink_inst.r_Count_2Z0Z_20 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_20 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_19 ;
    wire \led_blink_inst.r_Count_2Z0Z_21 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_20 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_21 ;
    wire \led_blink_inst.un2_r_Count_2_1_cry_22 ;
    wire \led_blink_inst.r_Count_2Z0Z_23 ;
    wire \led_blink_inst.o_LED_23_17 ;
    wire \led_blink_inst.o_LED_23_16 ;
    wire \led_blink_inst.r_Count_2_RNO_0Z0Z_22 ;
    wire \led_blink_inst.o_LED_23_21 ;
    wire \led_blink_inst.r_Count_2Z0Z_22 ;
    wire \led_blink_inst.o_LED_33_14 ;
    wire \led_blink_inst.o_LED_33_13 ;
    wire \led_blink_inst.o_LED_33_12_cascade_ ;
    wire \led_blink_inst.o_LED_33_21_cascade_ ;
    wire o_LED_3_c;
    wire \led_blink_inst.o_LED_33_16_cascade_ ;
    wire \led_blink_inst.o_LED_33_15 ;
    wire \led_blink_inst.o_LED_33_17 ;
    wire \led_blink_inst.o_LED_33_16 ;
    wire \led_blink_inst.o_LED_33_21 ;
    wire bfn_11_6_0_;
    wire \led_blink_inst.un2_r_Count_4_1_cry_1 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_2 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_3 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_4 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_5 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_6 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_7 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_8 ;
    wire bfn_11_7_0_;
    wire \led_blink_inst.un2_r_Count_4_1_cry_9 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_10 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_11 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_12 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_13 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_14 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_15 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_16 ;
    wire bfn_11_8_0_;
    wire \led_blink_inst.un2_r_Count_4_1_cry_17 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_18 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_19 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_20 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_21 ;
    wire \led_blink_inst.un2_r_Count_4_1_cry_22 ;
    wire \led_blink_inst.r_Count_3Z0Z_1 ;
    wire \led_blink_inst.r_Count_3Z0Z_0 ;
    wire bfn_12_3_0_;
    wire \led_blink_inst.r_Count_3Z0Z_2 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_1 ;
    wire \led_blink_inst.r_Count_3Z0Z_3 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_2 ;
    wire \led_blink_inst.r_Count_3Z0Z_4 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_3 ;
    wire \led_blink_inst.r_Count_3Z0Z_5 ;
    wire \led_blink_inst.r_Count_3_RNO_0Z0Z_5 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_4 ;
    wire \led_blink_inst.r_Count_3Z0Z_6 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_5 ;
    wire \led_blink_inst.r_Count_3Z0Z_7 ;
    wire \led_blink_inst.r_Count_3_RNO_0Z0Z_7 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_6 ;
    wire \led_blink_inst.r_Count_3Z0Z_8 ;
    wire \led_blink_inst.r_Count_3_RNO_0Z0Z_8 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_7 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_8 ;
    wire \led_blink_inst.r_Count_3Z0Z_9 ;
    wire bfn_12_4_0_;
    wire \led_blink_inst.r_Count_3Z0Z_10 ;
    wire \led_blink_inst.r_Count_3_RNO_0Z0Z_10 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_9 ;
    wire \led_blink_inst.r_Count_3Z0Z_11 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_10 ;
    wire \led_blink_inst.r_Count_3Z0Z_12 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_11 ;
    wire \led_blink_inst.r_Count_3Z0Z_13 ;
    wire \led_blink_inst.r_Count_3_RNO_0Z0Z_13 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_12 ;
    wire \led_blink_inst.r_Count_3Z0Z_14 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_13 ;
    wire \led_blink_inst.r_Count_3Z0Z_15 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_14 ;
    wire \led_blink_inst.r_Count_3Z0Z_16 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_15 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_16 ;
    wire \led_blink_inst.r_Count_3Z0Z_17 ;
    wire \led_blink_inst.r_Count_3_RNO_0Z0Z_17 ;
    wire bfn_12_5_0_;
    wire \led_blink_inst.r_Count_3Z0Z_18 ;
    wire \led_blink_inst.r_Count_3_RNO_0Z0Z_18 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_17 ;
    wire \led_blink_inst.r_Count_3Z0Z_19 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_18 ;
    wire \led_blink_inst.r_Count_3Z0Z_20 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_19 ;
    wire \led_blink_inst.r_Count_3Z0Z_21 ;
    wire \led_blink_inst.r_Count_3_RNO_0Z0Z_21 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_20 ;
    wire \led_blink_inst.r_Count_3Z0Z_22 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_21 ;
    wire \led_blink_inst.un2_r_Count_3_1_cry_22 ;
    wire \led_blink_inst.r_Count_3Z0Z_23 ;
    wire \led_blink_inst.r_Count_4_RNO_0Z0Z_4 ;
    wire \led_blink_inst.r_Count_4_RNO_0Z0Z_7 ;
    wire \led_blink_inst.r_Count_4_RNO_0Z0Z_6 ;
    wire \led_blink_inst.r_Count_4_RNO_0Z0Z_9 ;
    wire \led_blink_inst.r_Count_4Z0Z_6 ;
    wire \led_blink_inst.r_Count_4Z0Z_9 ;
    wire \led_blink_inst.r_Count_4Z0Z_7 ;
    wire \led_blink_inst.r_Count_4Z0Z_4 ;
    wire \led_blink_inst.r_Count_4Z0Z_8 ;
    wire \led_blink_inst.r_Count_4Z0Z_10 ;
    wire \led_blink_inst.r_Count_4Z0Z_13 ;
    wire \led_blink_inst.r_Count_4Z0Z_5 ;
    wire \led_blink_inst.o_LED_43_16_cascade_ ;
    wire \led_blink_inst.r_Count_4_RNO_0Z0Z_16 ;
    wire \led_blink_inst.r_Count_4_RNO_0Z0Z_12 ;
    wire \led_blink_inst.r_Count_4Z0Z_14 ;
    wire \led_blink_inst.r_Count_4Z0Z_23 ;
    wire \led_blink_inst.r_Count_4Z0Z_21 ;
    wire \led_blink_inst.r_Count_4Z0Z_3 ;
    wire \led_blink_inst.o_LED_43_12_cascade_ ;
    wire \led_blink_inst.o_LED_43_14 ;
    wire \led_blink_inst.r_Count_4Z0Z_11 ;
    wire \led_blink_inst.r_Count_4Z0Z_2 ;
    wire \led_blink_inst.r_Count_4Z0Z_18 ;
    wire \led_blink_inst.r_Count_4Z0Z_15 ;
    wire \led_blink_inst.o_LED_43_13 ;
    wire \led_blink_inst.r_Count_4Z0Z_19 ;
    wire \led_blink_inst.r_Count_4Z0Z_0 ;
    wire \led_blink_inst.r_Count_4Z0Z_22 ;
    wire \led_blink_inst.r_Count_4Z0Z_1 ;
    wire \led_blink_inst.o_LED_43_17_cascade_ ;
    wire o_LED_4_c;
    wire \led_blink_inst.r_Count_4_RNO_0Z0Z_20 ;
    wire \led_blink_inst.o_LED_43_17 ;
    wire \led_blink_inst.o_LED_43_16 ;
    wire \led_blink_inst.r_Count_4_RNO_0Z0Z_17 ;
    wire \led_blink_inst.o_LED_43_21 ;
    wire i_Clk_c_g;
    wire \led_blink_inst.r_Count_4Z0Z_12 ;
    wire \led_blink_inst.r_Count_4Z0Z_16 ;
    wire \led_blink_inst.r_Count_4Z0Z_17 ;
    wire \led_blink_inst.r_Count_4Z0Z_20 ;
    wire \led_blink_inst.o_LED_43_15 ;
    wire _gnd_net_;

    PRE_IO_GBUF i_Clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__5321),
            .GLOBALBUFFEROUTPUT(i_Clk_c_g));
    IO_PAD i_Clk_ibuf_gb_io_iopad (
            .OE(N__5323),
            .DIN(N__5322),
            .DOUT(N__5321),
            .PACKAGEPIN(i_Clk));
    defparam i_Clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam i_Clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Clk_ibuf_gb_io_preio (
            .PADOEN(N__5323),
            .PADOUT(N__5322),
            .PADIN(N__5321),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_1_obuf_iopad (
            .OE(N__5312),
            .DIN(N__5311),
            .DOUT(N__5310),
            .PACKAGEPIN(o_LED_1));
    defparam o_LED_1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_1_obuf_preio (
            .PADOEN(N__5312),
            .PADOUT(N__5311),
            .PADIN(N__5310),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2275),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_2_obuf_iopad (
            .OE(N__5303),
            .DIN(N__5302),
            .DOUT(N__5301),
            .PACKAGEPIN(o_LED_2));
    defparam o_LED_2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_2_obuf_preio (
            .PADOEN(N__5303),
            .PADOUT(N__5302),
            .PADIN(N__5301),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2824),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_3_obuf_iopad (
            .OE(N__5294),
            .DIN(N__5293),
            .DOUT(N__5292),
            .PACKAGEPIN(o_LED_3));
    defparam o_LED_3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_3_obuf_preio (
            .PADOEN(N__5294),
            .PADOUT(N__5293),
            .PADIN(N__5292),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3871),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_4_obuf_iopad (
            .OE(N__5285),
            .DIN(N__5284),
            .DOUT(N__5283),
            .PACKAGEPIN(o_LED_4));
    defparam o_LED_4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_4_obuf_preio (
            .PADOEN(N__5285),
            .PADOUT(N__5284),
            .PADIN(N__5283),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5110),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__1195 (
            .O(N__5266),
            .I(\led_blink_inst.o_LED_43_12_cascade_ ));
    InMux I__1194 (
            .O(N__5263),
            .I(N__5260));
    LocalMux I__1193 (
            .O(N__5260),
            .I(\led_blink_inst.o_LED_43_14 ));
    InMux I__1192 (
            .O(N__5257),
            .I(N__5253));
    InMux I__1191 (
            .O(N__5256),
            .I(N__5250));
    LocalMux I__1190 (
            .O(N__5253),
            .I(\led_blink_inst.r_Count_4Z0Z_11 ));
    LocalMux I__1189 (
            .O(N__5250),
            .I(\led_blink_inst.r_Count_4Z0Z_11 ));
    InMux I__1188 (
            .O(N__5245),
            .I(N__5241));
    InMux I__1187 (
            .O(N__5244),
            .I(N__5238));
    LocalMux I__1186 (
            .O(N__5241),
            .I(\led_blink_inst.r_Count_4Z0Z_2 ));
    LocalMux I__1185 (
            .O(N__5238),
            .I(\led_blink_inst.r_Count_4Z0Z_2 ));
    CascadeMux I__1184 (
            .O(N__5233),
            .I(N__5229));
    CascadeMux I__1183 (
            .O(N__5232),
            .I(N__5226));
    InMux I__1182 (
            .O(N__5229),
            .I(N__5223));
    InMux I__1181 (
            .O(N__5226),
            .I(N__5220));
    LocalMux I__1180 (
            .O(N__5223),
            .I(\led_blink_inst.r_Count_4Z0Z_18 ));
    LocalMux I__1179 (
            .O(N__5220),
            .I(\led_blink_inst.r_Count_4Z0Z_18 ));
    CascadeMux I__1178 (
            .O(N__5215),
            .I(N__5211));
    InMux I__1177 (
            .O(N__5214),
            .I(N__5208));
    InMux I__1176 (
            .O(N__5211),
            .I(N__5205));
    LocalMux I__1175 (
            .O(N__5208),
            .I(\led_blink_inst.r_Count_4Z0Z_15 ));
    LocalMux I__1174 (
            .O(N__5205),
            .I(\led_blink_inst.r_Count_4Z0Z_15 ));
    InMux I__1173 (
            .O(N__5200),
            .I(N__5197));
    LocalMux I__1172 (
            .O(N__5197),
            .I(N__5194));
    Odrv4 I__1171 (
            .O(N__5194),
            .I(\led_blink_inst.o_LED_43_13 ));
    CascadeMux I__1170 (
            .O(N__5191),
            .I(N__5187));
    InMux I__1169 (
            .O(N__5190),
            .I(N__5184));
    InMux I__1168 (
            .O(N__5187),
            .I(N__5181));
    LocalMux I__1167 (
            .O(N__5184),
            .I(\led_blink_inst.r_Count_4Z0Z_19 ));
    LocalMux I__1166 (
            .O(N__5181),
            .I(\led_blink_inst.r_Count_4Z0Z_19 ));
    InMux I__1165 (
            .O(N__5176),
            .I(N__5171));
    InMux I__1164 (
            .O(N__5175),
            .I(N__5165));
    InMux I__1163 (
            .O(N__5174),
            .I(N__5165));
    LocalMux I__1162 (
            .O(N__5171),
            .I(N__5162));
    InMux I__1161 (
            .O(N__5170),
            .I(N__5159));
    LocalMux I__1160 (
            .O(N__5165),
            .I(\led_blink_inst.r_Count_4Z0Z_0 ));
    Odrv4 I__1159 (
            .O(N__5162),
            .I(\led_blink_inst.r_Count_4Z0Z_0 ));
    LocalMux I__1158 (
            .O(N__5159),
            .I(\led_blink_inst.r_Count_4Z0Z_0 ));
    CascadeMux I__1157 (
            .O(N__5152),
            .I(N__5148));
    InMux I__1156 (
            .O(N__5151),
            .I(N__5145));
    InMux I__1155 (
            .O(N__5148),
            .I(N__5142));
    LocalMux I__1154 (
            .O(N__5145),
            .I(\led_blink_inst.r_Count_4Z0Z_22 ));
    LocalMux I__1153 (
            .O(N__5142),
            .I(\led_blink_inst.r_Count_4Z0Z_22 ));
    InMux I__1152 (
            .O(N__5137),
            .I(N__5132));
    CascadeMux I__1151 (
            .O(N__5136),
            .I(N__5129));
    InMux I__1150 (
            .O(N__5135),
            .I(N__5126));
    LocalMux I__1149 (
            .O(N__5132),
            .I(N__5123));
    InMux I__1148 (
            .O(N__5129),
            .I(N__5120));
    LocalMux I__1147 (
            .O(N__5126),
            .I(\led_blink_inst.r_Count_4Z0Z_1 ));
    Odrv4 I__1146 (
            .O(N__5123),
            .I(\led_blink_inst.r_Count_4Z0Z_1 ));
    LocalMux I__1145 (
            .O(N__5120),
            .I(\led_blink_inst.r_Count_4Z0Z_1 ));
    CascadeMux I__1144 (
            .O(N__5113),
            .I(\led_blink_inst.o_LED_43_17_cascade_ ));
    IoInMux I__1143 (
            .O(N__5110),
            .I(N__5106));
    InMux I__1142 (
            .O(N__5109),
            .I(N__5103));
    LocalMux I__1141 (
            .O(N__5106),
            .I(o_LED_4_c));
    LocalMux I__1140 (
            .O(N__5103),
            .I(o_LED_4_c));
    InMux I__1139 (
            .O(N__5098),
            .I(N__5095));
    LocalMux I__1138 (
            .O(N__5095),
            .I(\led_blink_inst.r_Count_4_RNO_0Z0Z_20 ));
    CascadeMux I__1137 (
            .O(N__5092),
            .I(N__5083));
    CascadeMux I__1136 (
            .O(N__5091),
            .I(N__5080));
    InMux I__1135 (
            .O(N__5090),
            .I(N__5073));
    InMux I__1134 (
            .O(N__5089),
            .I(N__5073));
    InMux I__1133 (
            .O(N__5088),
            .I(N__5062));
    InMux I__1132 (
            .O(N__5087),
            .I(N__5062));
    InMux I__1131 (
            .O(N__5086),
            .I(N__5062));
    InMux I__1130 (
            .O(N__5083),
            .I(N__5062));
    InMux I__1129 (
            .O(N__5080),
            .I(N__5062));
    InMux I__1128 (
            .O(N__5079),
            .I(N__5057));
    InMux I__1127 (
            .O(N__5078),
            .I(N__5057));
    LocalMux I__1126 (
            .O(N__5073),
            .I(N__5054));
    LocalMux I__1125 (
            .O(N__5062),
            .I(\led_blink_inst.o_LED_43_17 ));
    LocalMux I__1124 (
            .O(N__5057),
            .I(\led_blink_inst.o_LED_43_17 ));
    Odrv4 I__1123 (
            .O(N__5054),
            .I(\led_blink_inst.o_LED_43_17 ));
    InMux I__1122 (
            .O(N__5047),
            .I(N__5041));
    InMux I__1121 (
            .O(N__5046),
            .I(N__5041));
    LocalMux I__1120 (
            .O(N__5041),
            .I(N__5031));
    InMux I__1119 (
            .O(N__5040),
            .I(N__5022));
    InMux I__1118 (
            .O(N__5039),
            .I(N__5022));
    InMux I__1117 (
            .O(N__5038),
            .I(N__5022));
    InMux I__1116 (
            .O(N__5037),
            .I(N__5022));
    InMux I__1115 (
            .O(N__5036),
            .I(N__5015));
    InMux I__1114 (
            .O(N__5035),
            .I(N__5015));
    InMux I__1113 (
            .O(N__5034),
            .I(N__5015));
    Odrv4 I__1112 (
            .O(N__5031),
            .I(\led_blink_inst.o_LED_43_16 ));
    LocalMux I__1111 (
            .O(N__5022),
            .I(\led_blink_inst.o_LED_43_16 ));
    LocalMux I__1110 (
            .O(N__5015),
            .I(\led_blink_inst.o_LED_43_16 ));
    CascadeMux I__1109 (
            .O(N__5008),
            .I(N__5005));
    InMux I__1108 (
            .O(N__5005),
            .I(N__5002));
    LocalMux I__1107 (
            .O(N__5002),
            .I(\led_blink_inst.r_Count_4_RNO_0Z0Z_17 ));
    CascadeMux I__1106 (
            .O(N__4999),
            .I(N__4995));
    InMux I__1105 (
            .O(N__4998),
            .I(N__4984));
    InMux I__1104 (
            .O(N__4995),
            .I(N__4984));
    CascadeMux I__1103 (
            .O(N__4994),
            .I(N__4979));
    InMux I__1102 (
            .O(N__4993),
            .I(N__4968));
    InMux I__1101 (
            .O(N__4992),
            .I(N__4968));
    InMux I__1100 (
            .O(N__4991),
            .I(N__4968));
    InMux I__1099 (
            .O(N__4990),
            .I(N__4968));
    InMux I__1098 (
            .O(N__4989),
            .I(N__4968));
    LocalMux I__1097 (
            .O(N__4984),
            .I(N__4965));
    InMux I__1096 (
            .O(N__4983),
            .I(N__4958));
    InMux I__1095 (
            .O(N__4982),
            .I(N__4958));
    InMux I__1094 (
            .O(N__4979),
            .I(N__4958));
    LocalMux I__1093 (
            .O(N__4968),
            .I(\led_blink_inst.o_LED_43_21 ));
    Odrv4 I__1092 (
            .O(N__4965),
            .I(\led_blink_inst.o_LED_43_21 ));
    LocalMux I__1091 (
            .O(N__4958),
            .I(\led_blink_inst.o_LED_43_21 ));
    ClkMux I__1090 (
            .O(N__4951),
            .I(N__4876));
    ClkMux I__1089 (
            .O(N__4950),
            .I(N__4876));
    ClkMux I__1088 (
            .O(N__4949),
            .I(N__4876));
    ClkMux I__1087 (
            .O(N__4948),
            .I(N__4876));
    ClkMux I__1086 (
            .O(N__4947),
            .I(N__4876));
    ClkMux I__1085 (
            .O(N__4946),
            .I(N__4876));
    ClkMux I__1084 (
            .O(N__4945),
            .I(N__4876));
    ClkMux I__1083 (
            .O(N__4944),
            .I(N__4876));
    ClkMux I__1082 (
            .O(N__4943),
            .I(N__4876));
    ClkMux I__1081 (
            .O(N__4942),
            .I(N__4876));
    ClkMux I__1080 (
            .O(N__4941),
            .I(N__4876));
    ClkMux I__1079 (
            .O(N__4940),
            .I(N__4876));
    ClkMux I__1078 (
            .O(N__4939),
            .I(N__4876));
    ClkMux I__1077 (
            .O(N__4938),
            .I(N__4876));
    ClkMux I__1076 (
            .O(N__4937),
            .I(N__4876));
    ClkMux I__1075 (
            .O(N__4936),
            .I(N__4876));
    ClkMux I__1074 (
            .O(N__4935),
            .I(N__4876));
    ClkMux I__1073 (
            .O(N__4934),
            .I(N__4876));
    ClkMux I__1072 (
            .O(N__4933),
            .I(N__4876));
    ClkMux I__1071 (
            .O(N__4932),
            .I(N__4876));
    ClkMux I__1070 (
            .O(N__4931),
            .I(N__4876));
    ClkMux I__1069 (
            .O(N__4930),
            .I(N__4876));
    ClkMux I__1068 (
            .O(N__4929),
            .I(N__4876));
    ClkMux I__1067 (
            .O(N__4928),
            .I(N__4876));
    ClkMux I__1066 (
            .O(N__4927),
            .I(N__4876));
    GlobalMux I__1065 (
            .O(N__4876),
            .I(N__4873));
    gio2CtrlBuf I__1064 (
            .O(N__4873),
            .I(i_Clk_c_g));
    InMux I__1063 (
            .O(N__4870),
            .I(N__4866));
    InMux I__1062 (
            .O(N__4869),
            .I(N__4863));
    LocalMux I__1061 (
            .O(N__4866),
            .I(N__4860));
    LocalMux I__1060 (
            .O(N__4863),
            .I(\led_blink_inst.r_Count_4Z0Z_12 ));
    Odrv4 I__1059 (
            .O(N__4860),
            .I(\led_blink_inst.r_Count_4Z0Z_12 ));
    CascadeMux I__1058 (
            .O(N__4855),
            .I(N__4851));
    InMux I__1057 (
            .O(N__4854),
            .I(N__4848));
    InMux I__1056 (
            .O(N__4851),
            .I(N__4845));
    LocalMux I__1055 (
            .O(N__4848),
            .I(\led_blink_inst.r_Count_4Z0Z_16 ));
    LocalMux I__1054 (
            .O(N__4845),
            .I(\led_blink_inst.r_Count_4Z0Z_16 ));
    CascadeMux I__1053 (
            .O(N__4840),
            .I(N__4836));
    InMux I__1052 (
            .O(N__4839),
            .I(N__4833));
    InMux I__1051 (
            .O(N__4836),
            .I(N__4830));
    LocalMux I__1050 (
            .O(N__4833),
            .I(\led_blink_inst.r_Count_4Z0Z_17 ));
    LocalMux I__1049 (
            .O(N__4830),
            .I(\led_blink_inst.r_Count_4Z0Z_17 ));
    InMux I__1048 (
            .O(N__4825),
            .I(N__4821));
    InMux I__1047 (
            .O(N__4824),
            .I(N__4818));
    LocalMux I__1046 (
            .O(N__4821),
            .I(\led_blink_inst.r_Count_4Z0Z_20 ));
    LocalMux I__1045 (
            .O(N__4818),
            .I(\led_blink_inst.r_Count_4Z0Z_20 ));
    InMux I__1044 (
            .O(N__4813),
            .I(N__4810));
    LocalMux I__1043 (
            .O(N__4810),
            .I(\led_blink_inst.o_LED_43_15 ));
    InMux I__1042 (
            .O(N__4807),
            .I(N__4804));
    LocalMux I__1041 (
            .O(N__4804),
            .I(\led_blink_inst.r_Count_4_RNO_0Z0Z_9 ));
    InMux I__1040 (
            .O(N__4801),
            .I(N__4797));
    InMux I__1039 (
            .O(N__4800),
            .I(N__4794));
    LocalMux I__1038 (
            .O(N__4797),
            .I(\led_blink_inst.r_Count_4Z0Z_6 ));
    LocalMux I__1037 (
            .O(N__4794),
            .I(\led_blink_inst.r_Count_4Z0Z_6 ));
    InMux I__1036 (
            .O(N__4789),
            .I(N__4785));
    InMux I__1035 (
            .O(N__4788),
            .I(N__4782));
    LocalMux I__1034 (
            .O(N__4785),
            .I(\led_blink_inst.r_Count_4Z0Z_9 ));
    LocalMux I__1033 (
            .O(N__4782),
            .I(\led_blink_inst.r_Count_4Z0Z_9 ));
    CascadeMux I__1032 (
            .O(N__4777),
            .I(N__4774));
    InMux I__1031 (
            .O(N__4774),
            .I(N__4770));
    InMux I__1030 (
            .O(N__4773),
            .I(N__4767));
    LocalMux I__1029 (
            .O(N__4770),
            .I(\led_blink_inst.r_Count_4Z0Z_7 ));
    LocalMux I__1028 (
            .O(N__4767),
            .I(\led_blink_inst.r_Count_4Z0Z_7 ));
    InMux I__1027 (
            .O(N__4762),
            .I(N__4758));
    InMux I__1026 (
            .O(N__4761),
            .I(N__4755));
    LocalMux I__1025 (
            .O(N__4758),
            .I(\led_blink_inst.r_Count_4Z0Z_4 ));
    LocalMux I__1024 (
            .O(N__4755),
            .I(\led_blink_inst.r_Count_4Z0Z_4 ));
    CascadeMux I__1023 (
            .O(N__4750),
            .I(N__4746));
    InMux I__1022 (
            .O(N__4749),
            .I(N__4743));
    InMux I__1021 (
            .O(N__4746),
            .I(N__4740));
    LocalMux I__1020 (
            .O(N__4743),
            .I(\led_blink_inst.r_Count_4Z0Z_8 ));
    LocalMux I__1019 (
            .O(N__4740),
            .I(\led_blink_inst.r_Count_4Z0Z_8 ));
    InMux I__1018 (
            .O(N__4735),
            .I(N__4731));
    InMux I__1017 (
            .O(N__4734),
            .I(N__4728));
    LocalMux I__1016 (
            .O(N__4731),
            .I(\led_blink_inst.r_Count_4Z0Z_10 ));
    LocalMux I__1015 (
            .O(N__4728),
            .I(\led_blink_inst.r_Count_4Z0Z_10 ));
    CascadeMux I__1014 (
            .O(N__4723),
            .I(N__4719));
    CascadeMux I__1013 (
            .O(N__4722),
            .I(N__4716));
    InMux I__1012 (
            .O(N__4719),
            .I(N__4713));
    InMux I__1011 (
            .O(N__4716),
            .I(N__4710));
    LocalMux I__1010 (
            .O(N__4713),
            .I(\led_blink_inst.r_Count_4Z0Z_13 ));
    LocalMux I__1009 (
            .O(N__4710),
            .I(\led_blink_inst.r_Count_4Z0Z_13 ));
    CascadeMux I__1008 (
            .O(N__4705),
            .I(N__4701));
    InMux I__1007 (
            .O(N__4704),
            .I(N__4698));
    InMux I__1006 (
            .O(N__4701),
            .I(N__4695));
    LocalMux I__1005 (
            .O(N__4698),
            .I(\led_blink_inst.r_Count_4Z0Z_5 ));
    LocalMux I__1004 (
            .O(N__4695),
            .I(\led_blink_inst.r_Count_4Z0Z_5 ));
    CascadeMux I__1003 (
            .O(N__4690),
            .I(\led_blink_inst.o_LED_43_16_cascade_ ));
    InMux I__1002 (
            .O(N__4687),
            .I(N__4684));
    LocalMux I__1001 (
            .O(N__4684),
            .I(\led_blink_inst.r_Count_4_RNO_0Z0Z_16 ));
    CascadeMux I__1000 (
            .O(N__4681),
            .I(N__4678));
    InMux I__999 (
            .O(N__4678),
            .I(N__4675));
    LocalMux I__998 (
            .O(N__4675),
            .I(\led_blink_inst.r_Count_4_RNO_0Z0Z_12 ));
    InMux I__997 (
            .O(N__4672),
            .I(N__4669));
    LocalMux I__996 (
            .O(N__4669),
            .I(N__4665));
    InMux I__995 (
            .O(N__4668),
            .I(N__4662));
    Odrv4 I__994 (
            .O(N__4665),
            .I(\led_blink_inst.r_Count_4Z0Z_14 ));
    LocalMux I__993 (
            .O(N__4662),
            .I(\led_blink_inst.r_Count_4Z0Z_14 ));
    InMux I__992 (
            .O(N__4657),
            .I(N__4653));
    InMux I__991 (
            .O(N__4656),
            .I(N__4650));
    LocalMux I__990 (
            .O(N__4653),
            .I(\led_blink_inst.r_Count_4Z0Z_23 ));
    LocalMux I__989 (
            .O(N__4650),
            .I(\led_blink_inst.r_Count_4Z0Z_23 ));
    CascadeMux I__988 (
            .O(N__4645),
            .I(N__4641));
    InMux I__987 (
            .O(N__4644),
            .I(N__4638));
    InMux I__986 (
            .O(N__4641),
            .I(N__4635));
    LocalMux I__985 (
            .O(N__4638),
            .I(\led_blink_inst.r_Count_4Z0Z_21 ));
    LocalMux I__984 (
            .O(N__4635),
            .I(\led_blink_inst.r_Count_4Z0Z_21 ));
    InMux I__983 (
            .O(N__4630),
            .I(N__4626));
    InMux I__982 (
            .O(N__4629),
            .I(N__4623));
    LocalMux I__981 (
            .O(N__4626),
            .I(\led_blink_inst.r_Count_4Z0Z_3 ));
    LocalMux I__980 (
            .O(N__4623),
            .I(\led_blink_inst.r_Count_4Z0Z_3 ));
    CascadeMux I__979 (
            .O(N__4618),
            .I(N__4614));
    InMux I__978 (
            .O(N__4617),
            .I(N__4611));
    InMux I__977 (
            .O(N__4614),
            .I(N__4608));
    LocalMux I__976 (
            .O(N__4611),
            .I(\led_blink_inst.r_Count_3Z0Z_18 ));
    LocalMux I__975 (
            .O(N__4608),
            .I(\led_blink_inst.r_Count_3Z0Z_18 ));
    CascadeMux I__974 (
            .O(N__4603),
            .I(N__4600));
    InMux I__973 (
            .O(N__4600),
            .I(N__4597));
    LocalMux I__972 (
            .O(N__4597),
            .I(\led_blink_inst.r_Count_3_RNO_0Z0Z_18 ));
    InMux I__971 (
            .O(N__4594),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_17 ));
    CascadeMux I__970 (
            .O(N__4591),
            .I(N__4587));
    CascadeMux I__969 (
            .O(N__4590),
            .I(N__4584));
    InMux I__968 (
            .O(N__4587),
            .I(N__4581));
    InMux I__967 (
            .O(N__4584),
            .I(N__4578));
    LocalMux I__966 (
            .O(N__4581),
            .I(\led_blink_inst.r_Count_3Z0Z_19 ));
    LocalMux I__965 (
            .O(N__4578),
            .I(\led_blink_inst.r_Count_3Z0Z_19 ));
    InMux I__964 (
            .O(N__4573),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_18 ));
    CascadeMux I__963 (
            .O(N__4570),
            .I(N__4566));
    InMux I__962 (
            .O(N__4569),
            .I(N__4563));
    InMux I__961 (
            .O(N__4566),
            .I(N__4560));
    LocalMux I__960 (
            .O(N__4563),
            .I(\led_blink_inst.r_Count_3Z0Z_20 ));
    LocalMux I__959 (
            .O(N__4560),
            .I(\led_blink_inst.r_Count_3Z0Z_20 ));
    InMux I__958 (
            .O(N__4555),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_19 ));
    CascadeMux I__957 (
            .O(N__4552),
            .I(N__4548));
    InMux I__956 (
            .O(N__4551),
            .I(N__4545));
    InMux I__955 (
            .O(N__4548),
            .I(N__4542));
    LocalMux I__954 (
            .O(N__4545),
            .I(\led_blink_inst.r_Count_3Z0Z_21 ));
    LocalMux I__953 (
            .O(N__4542),
            .I(\led_blink_inst.r_Count_3Z0Z_21 ));
    InMux I__952 (
            .O(N__4537),
            .I(N__4534));
    LocalMux I__951 (
            .O(N__4534),
            .I(\led_blink_inst.r_Count_3_RNO_0Z0Z_21 ));
    InMux I__950 (
            .O(N__4531),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_20 ));
    CascadeMux I__949 (
            .O(N__4528),
            .I(N__4524));
    InMux I__948 (
            .O(N__4527),
            .I(N__4521));
    InMux I__947 (
            .O(N__4524),
            .I(N__4518));
    LocalMux I__946 (
            .O(N__4521),
            .I(\led_blink_inst.r_Count_3Z0Z_22 ));
    LocalMux I__945 (
            .O(N__4518),
            .I(\led_blink_inst.r_Count_3Z0Z_22 ));
    InMux I__944 (
            .O(N__4513),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_21 ));
    InMux I__943 (
            .O(N__4510),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_22 ));
    CascadeMux I__942 (
            .O(N__4507),
            .I(N__4504));
    InMux I__941 (
            .O(N__4504),
            .I(N__4500));
    InMux I__940 (
            .O(N__4503),
            .I(N__4497));
    LocalMux I__939 (
            .O(N__4500),
            .I(N__4494));
    LocalMux I__938 (
            .O(N__4497),
            .I(\led_blink_inst.r_Count_3Z0Z_23 ));
    Odrv4 I__937 (
            .O(N__4494),
            .I(\led_blink_inst.r_Count_3Z0Z_23 ));
    CascadeMux I__936 (
            .O(N__4489),
            .I(N__4486));
    InMux I__935 (
            .O(N__4486),
            .I(N__4483));
    LocalMux I__934 (
            .O(N__4483),
            .I(N__4480));
    Odrv4 I__933 (
            .O(N__4480),
            .I(\led_blink_inst.r_Count_4_RNO_0Z0Z_4 ));
    InMux I__932 (
            .O(N__4477),
            .I(N__4474));
    LocalMux I__931 (
            .O(N__4474),
            .I(\led_blink_inst.r_Count_4_RNO_0Z0Z_7 ));
    CascadeMux I__930 (
            .O(N__4471),
            .I(N__4468));
    InMux I__929 (
            .O(N__4468),
            .I(N__4465));
    LocalMux I__928 (
            .O(N__4465),
            .I(\led_blink_inst.r_Count_4_RNO_0Z0Z_6 ));
    CascadeMux I__927 (
            .O(N__4462),
            .I(N__4458));
    CascadeMux I__926 (
            .O(N__4461),
            .I(N__4455));
    InMux I__925 (
            .O(N__4458),
            .I(N__4452));
    InMux I__924 (
            .O(N__4455),
            .I(N__4449));
    LocalMux I__923 (
            .O(N__4452),
            .I(\led_blink_inst.r_Count_3Z0Z_10 ));
    LocalMux I__922 (
            .O(N__4449),
            .I(\led_blink_inst.r_Count_3Z0Z_10 ));
    InMux I__921 (
            .O(N__4444),
            .I(N__4441));
    LocalMux I__920 (
            .O(N__4441),
            .I(\led_blink_inst.r_Count_3_RNO_0Z0Z_10 ));
    InMux I__919 (
            .O(N__4438),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_9 ));
    CascadeMux I__918 (
            .O(N__4435),
            .I(N__4431));
    CascadeMux I__917 (
            .O(N__4434),
            .I(N__4428));
    InMux I__916 (
            .O(N__4431),
            .I(N__4425));
    InMux I__915 (
            .O(N__4428),
            .I(N__4422));
    LocalMux I__914 (
            .O(N__4425),
            .I(\led_blink_inst.r_Count_3Z0Z_11 ));
    LocalMux I__913 (
            .O(N__4422),
            .I(\led_blink_inst.r_Count_3Z0Z_11 ));
    InMux I__912 (
            .O(N__4417),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_10 ));
    CascadeMux I__911 (
            .O(N__4414),
            .I(N__4410));
    InMux I__910 (
            .O(N__4413),
            .I(N__4407));
    InMux I__909 (
            .O(N__4410),
            .I(N__4404));
    LocalMux I__908 (
            .O(N__4407),
            .I(\led_blink_inst.r_Count_3Z0Z_12 ));
    LocalMux I__907 (
            .O(N__4404),
            .I(\led_blink_inst.r_Count_3Z0Z_12 ));
    InMux I__906 (
            .O(N__4399),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_11 ));
    InMux I__905 (
            .O(N__4396),
            .I(N__4392));
    InMux I__904 (
            .O(N__4395),
            .I(N__4389));
    LocalMux I__903 (
            .O(N__4392),
            .I(\led_blink_inst.r_Count_3Z0Z_13 ));
    LocalMux I__902 (
            .O(N__4389),
            .I(\led_blink_inst.r_Count_3Z0Z_13 ));
    InMux I__901 (
            .O(N__4384),
            .I(N__4381));
    LocalMux I__900 (
            .O(N__4381),
            .I(\led_blink_inst.r_Count_3_RNO_0Z0Z_13 ));
    InMux I__899 (
            .O(N__4378),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_12 ));
    InMux I__898 (
            .O(N__4375),
            .I(N__4372));
    LocalMux I__897 (
            .O(N__4372),
            .I(N__4368));
    InMux I__896 (
            .O(N__4371),
            .I(N__4365));
    Odrv4 I__895 (
            .O(N__4368),
            .I(\led_blink_inst.r_Count_3Z0Z_14 ));
    LocalMux I__894 (
            .O(N__4365),
            .I(\led_blink_inst.r_Count_3Z0Z_14 ));
    InMux I__893 (
            .O(N__4360),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_13 ));
    CascadeMux I__892 (
            .O(N__4357),
            .I(N__4353));
    InMux I__891 (
            .O(N__4356),
            .I(N__4350));
    InMux I__890 (
            .O(N__4353),
            .I(N__4347));
    LocalMux I__889 (
            .O(N__4350),
            .I(\led_blink_inst.r_Count_3Z0Z_15 ));
    LocalMux I__888 (
            .O(N__4347),
            .I(\led_blink_inst.r_Count_3Z0Z_15 ));
    InMux I__887 (
            .O(N__4342),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_14 ));
    CascadeMux I__886 (
            .O(N__4339),
            .I(N__4335));
    InMux I__885 (
            .O(N__4338),
            .I(N__4332));
    InMux I__884 (
            .O(N__4335),
            .I(N__4329));
    LocalMux I__883 (
            .O(N__4332),
            .I(\led_blink_inst.r_Count_3Z0Z_16 ));
    LocalMux I__882 (
            .O(N__4329),
            .I(\led_blink_inst.r_Count_3Z0Z_16 ));
    InMux I__881 (
            .O(N__4324),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_15 ));
    InMux I__880 (
            .O(N__4321),
            .I(N__4317));
    InMux I__879 (
            .O(N__4320),
            .I(N__4314));
    LocalMux I__878 (
            .O(N__4317),
            .I(\led_blink_inst.r_Count_3Z0Z_17 ));
    LocalMux I__877 (
            .O(N__4314),
            .I(\led_blink_inst.r_Count_3Z0Z_17 ));
    CascadeMux I__876 (
            .O(N__4309),
            .I(N__4306));
    InMux I__875 (
            .O(N__4306),
            .I(N__4303));
    LocalMux I__874 (
            .O(N__4303),
            .I(\led_blink_inst.r_Count_3_RNO_0Z0Z_17 ));
    InMux I__873 (
            .O(N__4300),
            .I(bfn_12_5_0_));
    InMux I__872 (
            .O(N__4297),
            .I(N__4293));
    InMux I__871 (
            .O(N__4296),
            .I(N__4290));
    LocalMux I__870 (
            .O(N__4293),
            .I(\led_blink_inst.r_Count_3Z0Z_2 ));
    LocalMux I__869 (
            .O(N__4290),
            .I(\led_blink_inst.r_Count_3Z0Z_2 ));
    InMux I__868 (
            .O(N__4285),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_1 ));
    InMux I__867 (
            .O(N__4282),
            .I(N__4278));
    InMux I__866 (
            .O(N__4281),
            .I(N__4275));
    LocalMux I__865 (
            .O(N__4278),
            .I(\led_blink_inst.r_Count_3Z0Z_3 ));
    LocalMux I__864 (
            .O(N__4275),
            .I(\led_blink_inst.r_Count_3Z0Z_3 ));
    InMux I__863 (
            .O(N__4270),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_2 ));
    CascadeMux I__862 (
            .O(N__4267),
            .I(N__4263));
    InMux I__861 (
            .O(N__4266),
            .I(N__4260));
    InMux I__860 (
            .O(N__4263),
            .I(N__4257));
    LocalMux I__859 (
            .O(N__4260),
            .I(\led_blink_inst.r_Count_3Z0Z_4 ));
    LocalMux I__858 (
            .O(N__4257),
            .I(\led_blink_inst.r_Count_3Z0Z_4 ));
    InMux I__857 (
            .O(N__4252),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_3 ));
    InMux I__856 (
            .O(N__4249),
            .I(N__4245));
    InMux I__855 (
            .O(N__4248),
            .I(N__4242));
    LocalMux I__854 (
            .O(N__4245),
            .I(\led_blink_inst.r_Count_3Z0Z_5 ));
    LocalMux I__853 (
            .O(N__4242),
            .I(\led_blink_inst.r_Count_3Z0Z_5 ));
    InMux I__852 (
            .O(N__4237),
            .I(N__4234));
    LocalMux I__851 (
            .O(N__4234),
            .I(\led_blink_inst.r_Count_3_RNO_0Z0Z_5 ));
    InMux I__850 (
            .O(N__4231),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_4 ));
    InMux I__849 (
            .O(N__4228),
            .I(N__4225));
    LocalMux I__848 (
            .O(N__4225),
            .I(N__4221));
    InMux I__847 (
            .O(N__4224),
            .I(N__4218));
    Odrv4 I__846 (
            .O(N__4221),
            .I(\led_blink_inst.r_Count_3Z0Z_6 ));
    LocalMux I__845 (
            .O(N__4218),
            .I(\led_blink_inst.r_Count_3Z0Z_6 ));
    InMux I__844 (
            .O(N__4213),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_5 ));
    InMux I__843 (
            .O(N__4210),
            .I(N__4207));
    LocalMux I__842 (
            .O(N__4207),
            .I(N__4203));
    InMux I__841 (
            .O(N__4206),
            .I(N__4200));
    Odrv4 I__840 (
            .O(N__4203),
            .I(\led_blink_inst.r_Count_3Z0Z_7 ));
    LocalMux I__839 (
            .O(N__4200),
            .I(\led_blink_inst.r_Count_3Z0Z_7 ));
    InMux I__838 (
            .O(N__4195),
            .I(N__4192));
    LocalMux I__837 (
            .O(N__4192),
            .I(\led_blink_inst.r_Count_3_RNO_0Z0Z_7 ));
    InMux I__836 (
            .O(N__4189),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_6 ));
    CascadeMux I__835 (
            .O(N__4186),
            .I(N__4182));
    InMux I__834 (
            .O(N__4185),
            .I(N__4179));
    InMux I__833 (
            .O(N__4182),
            .I(N__4176));
    LocalMux I__832 (
            .O(N__4179),
            .I(\led_blink_inst.r_Count_3Z0Z_8 ));
    LocalMux I__831 (
            .O(N__4176),
            .I(\led_blink_inst.r_Count_3Z0Z_8 ));
    CascadeMux I__830 (
            .O(N__4171),
            .I(N__4168));
    InMux I__829 (
            .O(N__4168),
            .I(N__4165));
    LocalMux I__828 (
            .O(N__4165),
            .I(N__4162));
    Odrv4 I__827 (
            .O(N__4162),
            .I(\led_blink_inst.r_Count_3_RNO_0Z0Z_8 ));
    InMux I__826 (
            .O(N__4159),
            .I(\led_blink_inst.un2_r_Count_3_1_cry_7 ));
    CascadeMux I__825 (
            .O(N__4156),
            .I(N__4152));
    InMux I__824 (
            .O(N__4155),
            .I(N__4149));
    InMux I__823 (
            .O(N__4152),
            .I(N__4146));
    LocalMux I__822 (
            .O(N__4149),
            .I(\led_blink_inst.r_Count_3Z0Z_9 ));
    LocalMux I__821 (
            .O(N__4146),
            .I(\led_blink_inst.r_Count_3Z0Z_9 ));
    InMux I__820 (
            .O(N__4141),
            .I(bfn_12_4_0_));
    InMux I__819 (
            .O(N__4138),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_15 ));
    InMux I__818 (
            .O(N__4135),
            .I(bfn_11_8_0_));
    InMux I__817 (
            .O(N__4132),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_17 ));
    InMux I__816 (
            .O(N__4129),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_18 ));
    InMux I__815 (
            .O(N__4126),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_19 ));
    InMux I__814 (
            .O(N__4123),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_20 ));
    InMux I__813 (
            .O(N__4120),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_21 ));
    InMux I__812 (
            .O(N__4117),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_22 ));
    InMux I__811 (
            .O(N__4114),
            .I(N__4107));
    InMux I__810 (
            .O(N__4113),
            .I(N__4107));
    InMux I__809 (
            .O(N__4112),
            .I(N__4104));
    LocalMux I__808 (
            .O(N__4107),
            .I(\led_blink_inst.r_Count_3Z0Z_1 ));
    LocalMux I__807 (
            .O(N__4104),
            .I(\led_blink_inst.r_Count_3Z0Z_1 ));
    CascadeMux I__806 (
            .O(N__4099),
            .I(N__4093));
    InMux I__805 (
            .O(N__4098),
            .I(N__4090));
    InMux I__804 (
            .O(N__4097),
            .I(N__4085));
    InMux I__803 (
            .O(N__4096),
            .I(N__4085));
    InMux I__802 (
            .O(N__4093),
            .I(N__4082));
    LocalMux I__801 (
            .O(N__4090),
            .I(\led_blink_inst.r_Count_3Z0Z_0 ));
    LocalMux I__800 (
            .O(N__4085),
            .I(\led_blink_inst.r_Count_3Z0Z_0 ));
    LocalMux I__799 (
            .O(N__4082),
            .I(\led_blink_inst.r_Count_3Z0Z_0 ));
    InMux I__798 (
            .O(N__4075),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_6 ));
    InMux I__797 (
            .O(N__4072),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_7 ));
    InMux I__796 (
            .O(N__4069),
            .I(bfn_11_7_0_));
    InMux I__795 (
            .O(N__4066),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_9 ));
    InMux I__794 (
            .O(N__4063),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_10 ));
    InMux I__793 (
            .O(N__4060),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_11 ));
    InMux I__792 (
            .O(N__4057),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_12 ));
    InMux I__791 (
            .O(N__4054),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_13 ));
    InMux I__790 (
            .O(N__4051),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_14 ));
    InMux I__789 (
            .O(N__4048),
            .I(N__4045));
    LocalMux I__788 (
            .O(N__4045),
            .I(\led_blink_inst.o_LED_33_15 ));
    InMux I__787 (
            .O(N__4042),
            .I(N__4029));
    InMux I__786 (
            .O(N__4041),
            .I(N__4029));
    InMux I__785 (
            .O(N__4040),
            .I(N__4029));
    CascadeMux I__784 (
            .O(N__4039),
            .I(N__4024));
    InMux I__783 (
            .O(N__4038),
            .I(N__4016));
    InMux I__782 (
            .O(N__4037),
            .I(N__4016));
    InMux I__781 (
            .O(N__4036),
            .I(N__4016));
    LocalMux I__780 (
            .O(N__4029),
            .I(N__4013));
    InMux I__779 (
            .O(N__4028),
            .I(N__4006));
    InMux I__778 (
            .O(N__4027),
            .I(N__4006));
    InMux I__777 (
            .O(N__4024),
            .I(N__4006));
    InMux I__776 (
            .O(N__4023),
            .I(N__4003));
    LocalMux I__775 (
            .O(N__4016),
            .I(\led_blink_inst.o_LED_33_17 ));
    Odrv4 I__774 (
            .O(N__4013),
            .I(\led_blink_inst.o_LED_33_17 ));
    LocalMux I__773 (
            .O(N__4006),
            .I(\led_blink_inst.o_LED_33_17 ));
    LocalMux I__772 (
            .O(N__4003),
            .I(\led_blink_inst.o_LED_33_17 ));
    InMux I__771 (
            .O(N__3994),
            .I(N__3979));
    InMux I__770 (
            .O(N__3993),
            .I(N__3979));
    InMux I__769 (
            .O(N__3992),
            .I(N__3979));
    InMux I__768 (
            .O(N__3991),
            .I(N__3972));
    InMux I__767 (
            .O(N__3990),
            .I(N__3972));
    InMux I__766 (
            .O(N__3989),
            .I(N__3972));
    InMux I__765 (
            .O(N__3988),
            .I(N__3965));
    InMux I__764 (
            .O(N__3987),
            .I(N__3965));
    InMux I__763 (
            .O(N__3986),
            .I(N__3965));
    LocalMux I__762 (
            .O(N__3979),
            .I(\led_blink_inst.o_LED_33_16 ));
    LocalMux I__761 (
            .O(N__3972),
            .I(\led_blink_inst.o_LED_33_16 ));
    LocalMux I__760 (
            .O(N__3965),
            .I(\led_blink_inst.o_LED_33_16 ));
    CascadeMux I__759 (
            .O(N__3958),
            .I(N__3951));
    CascadeMux I__758 (
            .O(N__3957),
            .I(N__3948));
    CascadeMux I__757 (
            .O(N__3956),
            .I(N__3943));
    CascadeMux I__756 (
            .O(N__3955),
            .I(N__3938));
    InMux I__755 (
            .O(N__3954),
            .I(N__3935));
    InMux I__754 (
            .O(N__3951),
            .I(N__3930));
    InMux I__753 (
            .O(N__3948),
            .I(N__3930));
    InMux I__752 (
            .O(N__3947),
            .I(N__3923));
    InMux I__751 (
            .O(N__3946),
            .I(N__3923));
    InMux I__750 (
            .O(N__3943),
            .I(N__3923));
    InMux I__749 (
            .O(N__3942),
            .I(N__3916));
    InMux I__748 (
            .O(N__3941),
            .I(N__3916));
    InMux I__747 (
            .O(N__3938),
            .I(N__3916));
    LocalMux I__746 (
            .O(N__3935),
            .I(\led_blink_inst.o_LED_33_21 ));
    LocalMux I__745 (
            .O(N__3930),
            .I(\led_blink_inst.o_LED_33_21 ));
    LocalMux I__744 (
            .O(N__3923),
            .I(\led_blink_inst.o_LED_33_21 ));
    LocalMux I__743 (
            .O(N__3916),
            .I(\led_blink_inst.o_LED_33_21 ));
    InMux I__742 (
            .O(N__3907),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_1 ));
    InMux I__741 (
            .O(N__3904),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_2 ));
    InMux I__740 (
            .O(N__3901),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_3 ));
    InMux I__739 (
            .O(N__3898),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_4 ));
    InMux I__738 (
            .O(N__3895),
            .I(\led_blink_inst.un2_r_Count_4_1_cry_5 ));
    InMux I__737 (
            .O(N__3892),
            .I(N__3889));
    LocalMux I__736 (
            .O(N__3889),
            .I(N__3886));
    Odrv4 I__735 (
            .O(N__3886),
            .I(\led_blink_inst.o_LED_33_14 ));
    InMux I__734 (
            .O(N__3883),
            .I(N__3880));
    LocalMux I__733 (
            .O(N__3880),
            .I(\led_blink_inst.o_LED_33_13 ));
    CascadeMux I__732 (
            .O(N__3877),
            .I(\led_blink_inst.o_LED_33_12_cascade_ ));
    CascadeMux I__731 (
            .O(N__3874),
            .I(\led_blink_inst.o_LED_33_21_cascade_ ));
    IoInMux I__730 (
            .O(N__3871),
            .I(N__3868));
    LocalMux I__729 (
            .O(N__3868),
            .I(N__3864));
    InMux I__728 (
            .O(N__3867),
            .I(N__3861));
    Span4Mux_s1_h I__727 (
            .O(N__3864),
            .I(N__3858));
    LocalMux I__726 (
            .O(N__3861),
            .I(N__3855));
    Odrv4 I__725 (
            .O(N__3858),
            .I(o_LED_3_c));
    Odrv4 I__724 (
            .O(N__3855),
            .I(o_LED_3_c));
    CascadeMux I__723 (
            .O(N__3850),
            .I(\led_blink_inst.o_LED_33_16_cascade_ ));
    CascadeMux I__722 (
            .O(N__3847),
            .I(N__3844));
    InMux I__721 (
            .O(N__3844),
            .I(N__3840));
    CascadeMux I__720 (
            .O(N__3843),
            .I(N__3837));
    LocalMux I__719 (
            .O(N__3840),
            .I(N__3834));
    InMux I__718 (
            .O(N__3837),
            .I(N__3831));
    Odrv4 I__717 (
            .O(N__3834),
            .I(\led_blink_inst.r_Count_2Z0Z_21 ));
    LocalMux I__716 (
            .O(N__3831),
            .I(\led_blink_inst.r_Count_2Z0Z_21 ));
    InMux I__715 (
            .O(N__3826),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_20 ));
    InMux I__714 (
            .O(N__3823),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_21 ));
    InMux I__713 (
            .O(N__3820),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_22 ));
    InMux I__712 (
            .O(N__3817),
            .I(N__3813));
    InMux I__711 (
            .O(N__3816),
            .I(N__3810));
    LocalMux I__710 (
            .O(N__3813),
            .I(N__3807));
    LocalMux I__709 (
            .O(N__3810),
            .I(\led_blink_inst.r_Count_2Z0Z_23 ));
    Odrv12 I__708 (
            .O(N__3807),
            .I(\led_blink_inst.r_Count_2Z0Z_23 ));
    InMux I__707 (
            .O(N__3802),
            .I(N__3798));
    CascadeMux I__706 (
            .O(N__3801),
            .I(N__3783));
    LocalMux I__705 (
            .O(N__3798),
            .I(N__3780));
    InMux I__704 (
            .O(N__3797),
            .I(N__3767));
    InMux I__703 (
            .O(N__3796),
            .I(N__3767));
    InMux I__702 (
            .O(N__3795),
            .I(N__3767));
    InMux I__701 (
            .O(N__3794),
            .I(N__3767));
    InMux I__700 (
            .O(N__3793),
            .I(N__3767));
    InMux I__699 (
            .O(N__3792),
            .I(N__3767));
    InMux I__698 (
            .O(N__3791),
            .I(N__3764));
    InMux I__697 (
            .O(N__3790),
            .I(N__3757));
    InMux I__696 (
            .O(N__3789),
            .I(N__3757));
    InMux I__695 (
            .O(N__3788),
            .I(N__3757));
    InMux I__694 (
            .O(N__3787),
            .I(N__3750));
    InMux I__693 (
            .O(N__3786),
            .I(N__3750));
    InMux I__692 (
            .O(N__3783),
            .I(N__3750));
    Odrv12 I__691 (
            .O(N__3780),
            .I(\led_blink_inst.o_LED_23_17 ));
    LocalMux I__690 (
            .O(N__3767),
            .I(\led_blink_inst.o_LED_23_17 ));
    LocalMux I__689 (
            .O(N__3764),
            .I(\led_blink_inst.o_LED_23_17 ));
    LocalMux I__688 (
            .O(N__3757),
            .I(\led_blink_inst.o_LED_23_17 ));
    LocalMux I__687 (
            .O(N__3750),
            .I(\led_blink_inst.o_LED_23_17 ));
    InMux I__686 (
            .O(N__3739),
            .I(N__3736));
    LocalMux I__685 (
            .O(N__3736),
            .I(N__3733));
    Span4Mux_v I__684 (
            .O(N__3733),
            .I(N__3718));
    InMux I__683 (
            .O(N__3732),
            .I(N__3705));
    InMux I__682 (
            .O(N__3731),
            .I(N__3705));
    InMux I__681 (
            .O(N__3730),
            .I(N__3705));
    InMux I__680 (
            .O(N__3729),
            .I(N__3705));
    InMux I__679 (
            .O(N__3728),
            .I(N__3705));
    InMux I__678 (
            .O(N__3727),
            .I(N__3705));
    InMux I__677 (
            .O(N__3726),
            .I(N__3698));
    InMux I__676 (
            .O(N__3725),
            .I(N__3698));
    InMux I__675 (
            .O(N__3724),
            .I(N__3698));
    InMux I__674 (
            .O(N__3723),
            .I(N__3691));
    InMux I__673 (
            .O(N__3722),
            .I(N__3691));
    InMux I__672 (
            .O(N__3721),
            .I(N__3691));
    Odrv4 I__671 (
            .O(N__3718),
            .I(\led_blink_inst.o_LED_23_16 ));
    LocalMux I__670 (
            .O(N__3705),
            .I(\led_blink_inst.o_LED_23_16 ));
    LocalMux I__669 (
            .O(N__3698),
            .I(\led_blink_inst.o_LED_23_16 ));
    LocalMux I__668 (
            .O(N__3691),
            .I(\led_blink_inst.o_LED_23_16 ));
    CascadeMux I__667 (
            .O(N__3682),
            .I(N__3679));
    InMux I__666 (
            .O(N__3679),
            .I(N__3676));
    LocalMux I__665 (
            .O(N__3676),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_22 ));
    InMux I__664 (
            .O(N__3673),
            .I(N__3666));
    CascadeMux I__663 (
            .O(N__3672),
            .I(N__3661));
    CascadeMux I__662 (
            .O(N__3671),
            .I(N__3657));
    CascadeMux I__661 (
            .O(N__3670),
            .I(N__3652));
    CascadeMux I__660 (
            .O(N__3669),
            .I(N__3647));
    LocalMux I__659 (
            .O(N__3666),
            .I(N__3643));
    InMux I__658 (
            .O(N__3665),
            .I(N__3630));
    InMux I__657 (
            .O(N__3664),
            .I(N__3630));
    InMux I__656 (
            .O(N__3661),
            .I(N__3630));
    InMux I__655 (
            .O(N__3660),
            .I(N__3630));
    InMux I__654 (
            .O(N__3657),
            .I(N__3630));
    InMux I__653 (
            .O(N__3656),
            .I(N__3630));
    InMux I__652 (
            .O(N__3655),
            .I(N__3627));
    InMux I__651 (
            .O(N__3652),
            .I(N__3620));
    InMux I__650 (
            .O(N__3651),
            .I(N__3620));
    InMux I__649 (
            .O(N__3650),
            .I(N__3620));
    InMux I__648 (
            .O(N__3647),
            .I(N__3615));
    InMux I__647 (
            .O(N__3646),
            .I(N__3615));
    Odrv4 I__646 (
            .O(N__3643),
            .I(\led_blink_inst.o_LED_23_21 ));
    LocalMux I__645 (
            .O(N__3630),
            .I(\led_blink_inst.o_LED_23_21 ));
    LocalMux I__644 (
            .O(N__3627),
            .I(\led_blink_inst.o_LED_23_21 ));
    LocalMux I__643 (
            .O(N__3620),
            .I(\led_blink_inst.o_LED_23_21 ));
    LocalMux I__642 (
            .O(N__3615),
            .I(\led_blink_inst.o_LED_23_21 ));
    CascadeMux I__641 (
            .O(N__3604),
            .I(N__3601));
    InMux I__640 (
            .O(N__3601),
            .I(N__3598));
    LocalMux I__639 (
            .O(N__3598),
            .I(N__3595));
    Span4Mux_h I__638 (
            .O(N__3595),
            .I(N__3591));
    InMux I__637 (
            .O(N__3594),
            .I(N__3588));
    Odrv4 I__636 (
            .O(N__3591),
            .I(\led_blink_inst.r_Count_2Z0Z_22 ));
    LocalMux I__635 (
            .O(N__3588),
            .I(\led_blink_inst.r_Count_2Z0Z_22 ));
    CascadeMux I__634 (
            .O(N__3583),
            .I(N__3580));
    InMux I__633 (
            .O(N__3580),
            .I(N__3577));
    LocalMux I__632 (
            .O(N__3577),
            .I(N__3573));
    InMux I__631 (
            .O(N__3576),
            .I(N__3570));
    Odrv12 I__630 (
            .O(N__3573),
            .I(\led_blink_inst.r_Count_2Z0Z_13 ));
    LocalMux I__629 (
            .O(N__3570),
            .I(\led_blink_inst.r_Count_2Z0Z_13 ));
    InMux I__628 (
            .O(N__3565),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_12 ));
    InMux I__627 (
            .O(N__3562),
            .I(N__3558));
    InMux I__626 (
            .O(N__3561),
            .I(N__3555));
    LocalMux I__625 (
            .O(N__3558),
            .I(\led_blink_inst.r_Count_2Z0Z_14 ));
    LocalMux I__624 (
            .O(N__3555),
            .I(\led_blink_inst.r_Count_2Z0Z_14 ));
    InMux I__623 (
            .O(N__3550),
            .I(N__3547));
    LocalMux I__622 (
            .O(N__3547),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_14 ));
    InMux I__621 (
            .O(N__3544),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_13 ));
    InMux I__620 (
            .O(N__3541),
            .I(N__3537));
    CascadeMux I__619 (
            .O(N__3540),
            .I(N__3534));
    LocalMux I__618 (
            .O(N__3537),
            .I(N__3531));
    InMux I__617 (
            .O(N__3534),
            .I(N__3528));
    Odrv4 I__616 (
            .O(N__3531),
            .I(\led_blink_inst.r_Count_2Z0Z_15 ));
    LocalMux I__615 (
            .O(N__3528),
            .I(\led_blink_inst.r_Count_2Z0Z_15 ));
    InMux I__614 (
            .O(N__3523),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_14 ));
    InMux I__613 (
            .O(N__3520),
            .I(N__3516));
    InMux I__612 (
            .O(N__3519),
            .I(N__3513));
    LocalMux I__611 (
            .O(N__3516),
            .I(N__3510));
    LocalMux I__610 (
            .O(N__3513),
            .I(\led_blink_inst.r_Count_2Z0Z_16 ));
    Odrv12 I__609 (
            .O(N__3510),
            .I(\led_blink_inst.r_Count_2Z0Z_16 ));
    InMux I__608 (
            .O(N__3505),
            .I(N__3502));
    LocalMux I__607 (
            .O(N__3502),
            .I(N__3499));
    Odrv12 I__606 (
            .O(N__3499),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_16 ));
    InMux I__605 (
            .O(N__3496),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_15 ));
    CascadeMux I__604 (
            .O(N__3493),
            .I(N__3490));
    InMux I__603 (
            .O(N__3490),
            .I(N__3486));
    InMux I__602 (
            .O(N__3489),
            .I(N__3483));
    LocalMux I__601 (
            .O(N__3486),
            .I(N__3480));
    LocalMux I__600 (
            .O(N__3483),
            .I(\led_blink_inst.r_Count_2Z0Z_17 ));
    Odrv4 I__599 (
            .O(N__3480),
            .I(\led_blink_inst.r_Count_2Z0Z_17 ));
    CascadeMux I__598 (
            .O(N__3475),
            .I(N__3472));
    InMux I__597 (
            .O(N__3472),
            .I(N__3469));
    LocalMux I__596 (
            .O(N__3469),
            .I(N__3466));
    Span4Mux_h I__595 (
            .O(N__3466),
            .I(N__3463));
    Odrv4 I__594 (
            .O(N__3463),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_17 ));
    InMux I__593 (
            .O(N__3460),
            .I(bfn_9_8_0_));
    CascadeMux I__592 (
            .O(N__3457),
            .I(N__3454));
    InMux I__591 (
            .O(N__3454),
            .I(N__3450));
    InMux I__590 (
            .O(N__3453),
            .I(N__3447));
    LocalMux I__589 (
            .O(N__3450),
            .I(N__3444));
    LocalMux I__588 (
            .O(N__3447),
            .I(\led_blink_inst.r_Count_2Z0Z_18 ));
    Odrv4 I__587 (
            .O(N__3444),
            .I(\led_blink_inst.r_Count_2Z0Z_18 ));
    InMux I__586 (
            .O(N__3439),
            .I(N__3436));
    LocalMux I__585 (
            .O(N__3436),
            .I(N__3433));
    Odrv4 I__584 (
            .O(N__3433),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_18 ));
    InMux I__583 (
            .O(N__3430),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_17 ));
    InMux I__582 (
            .O(N__3427),
            .I(N__3423));
    InMux I__581 (
            .O(N__3426),
            .I(N__3420));
    LocalMux I__580 (
            .O(N__3423),
            .I(N__3417));
    LocalMux I__579 (
            .O(N__3420),
            .I(\led_blink_inst.r_Count_2Z0Z_19 ));
    Odrv4 I__578 (
            .O(N__3417),
            .I(\led_blink_inst.r_Count_2Z0Z_19 ));
    CascadeMux I__577 (
            .O(N__3412),
            .I(N__3409));
    InMux I__576 (
            .O(N__3409),
            .I(N__3406));
    LocalMux I__575 (
            .O(N__3406),
            .I(N__3403));
    Odrv4 I__574 (
            .O(N__3403),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_19 ));
    InMux I__573 (
            .O(N__3400),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_18 ));
    CascadeMux I__572 (
            .O(N__3397),
            .I(N__3394));
    InMux I__571 (
            .O(N__3394),
            .I(N__3390));
    InMux I__570 (
            .O(N__3393),
            .I(N__3387));
    LocalMux I__569 (
            .O(N__3390),
            .I(N__3384));
    LocalMux I__568 (
            .O(N__3387),
            .I(\led_blink_inst.r_Count_2Z0Z_20 ));
    Odrv4 I__567 (
            .O(N__3384),
            .I(\led_blink_inst.r_Count_2Z0Z_20 ));
    CascadeMux I__566 (
            .O(N__3379),
            .I(N__3376));
    InMux I__565 (
            .O(N__3376),
            .I(N__3373));
    LocalMux I__564 (
            .O(N__3373),
            .I(N__3370));
    Odrv4 I__563 (
            .O(N__3370),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_20 ));
    InMux I__562 (
            .O(N__3367),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_19 ));
    InMux I__561 (
            .O(N__3364),
            .I(N__3360));
    InMux I__560 (
            .O(N__3363),
            .I(N__3357));
    LocalMux I__559 (
            .O(N__3360),
            .I(\led_blink_inst.r_Count_2Z0Z_5 ));
    LocalMux I__558 (
            .O(N__3357),
            .I(\led_blink_inst.r_Count_2Z0Z_5 ));
    InMux I__557 (
            .O(N__3352),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_4 ));
    InMux I__556 (
            .O(N__3349),
            .I(N__3345));
    InMux I__555 (
            .O(N__3348),
            .I(N__3342));
    LocalMux I__554 (
            .O(N__3345),
            .I(\led_blink_inst.r_Count_2Z0Z_6 ));
    LocalMux I__553 (
            .O(N__3342),
            .I(\led_blink_inst.r_Count_2Z0Z_6 ));
    InMux I__552 (
            .O(N__3337),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_5 ));
    CascadeMux I__551 (
            .O(N__3334),
            .I(N__3330));
    InMux I__550 (
            .O(N__3333),
            .I(N__3327));
    InMux I__549 (
            .O(N__3330),
            .I(N__3324));
    LocalMux I__548 (
            .O(N__3327),
            .I(\led_blink_inst.r_Count_2Z0Z_7 ));
    LocalMux I__547 (
            .O(N__3324),
            .I(\led_blink_inst.r_Count_2Z0Z_7 ));
    InMux I__546 (
            .O(N__3319),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_6 ));
    InMux I__545 (
            .O(N__3316),
            .I(N__3312));
    InMux I__544 (
            .O(N__3315),
            .I(N__3309));
    LocalMux I__543 (
            .O(N__3312),
            .I(\led_blink_inst.r_Count_2Z0Z_8 ));
    LocalMux I__542 (
            .O(N__3309),
            .I(\led_blink_inst.r_Count_2Z0Z_8 ));
    InMux I__541 (
            .O(N__3304),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_7 ));
    InMux I__540 (
            .O(N__3301),
            .I(N__3297));
    InMux I__539 (
            .O(N__3300),
            .I(N__3294));
    LocalMux I__538 (
            .O(N__3297),
            .I(N__3291));
    LocalMux I__537 (
            .O(N__3294),
            .I(N__3288));
    Odrv4 I__536 (
            .O(N__3291),
            .I(\led_blink_inst.r_Count_2Z0Z_9 ));
    Odrv4 I__535 (
            .O(N__3288),
            .I(\led_blink_inst.r_Count_2Z0Z_9 ));
    InMux I__534 (
            .O(N__3283),
            .I(N__3280));
    LocalMux I__533 (
            .O(N__3280),
            .I(N__3277));
    Odrv4 I__532 (
            .O(N__3277),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_9 ));
    InMux I__531 (
            .O(N__3274),
            .I(bfn_9_7_0_));
    CascadeMux I__530 (
            .O(N__3271),
            .I(N__3267));
    InMux I__529 (
            .O(N__3270),
            .I(N__3264));
    InMux I__528 (
            .O(N__3267),
            .I(N__3261));
    LocalMux I__527 (
            .O(N__3264),
            .I(\led_blink_inst.r_Count_2Z0Z_10 ));
    LocalMux I__526 (
            .O(N__3261),
            .I(\led_blink_inst.r_Count_2Z0Z_10 ));
    CascadeMux I__525 (
            .O(N__3256),
            .I(N__3253));
    InMux I__524 (
            .O(N__3253),
            .I(N__3250));
    LocalMux I__523 (
            .O(N__3250),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_10 ));
    InMux I__522 (
            .O(N__3247),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_9 ));
    CascadeMux I__521 (
            .O(N__3244),
            .I(N__3240));
    InMux I__520 (
            .O(N__3243),
            .I(N__3237));
    InMux I__519 (
            .O(N__3240),
            .I(N__3234));
    LocalMux I__518 (
            .O(N__3237),
            .I(N__3231));
    LocalMux I__517 (
            .O(N__3234),
            .I(\led_blink_inst.r_Count_2Z0Z_11 ));
    Odrv4 I__516 (
            .O(N__3231),
            .I(\led_blink_inst.r_Count_2Z0Z_11 ));
    CascadeMux I__515 (
            .O(N__3226),
            .I(N__3223));
    InMux I__514 (
            .O(N__3223),
            .I(N__3220));
    LocalMux I__513 (
            .O(N__3220),
            .I(N__3217));
    Odrv4 I__512 (
            .O(N__3217),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_11 ));
    InMux I__511 (
            .O(N__3214),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_10 ));
    CascadeMux I__510 (
            .O(N__3211),
            .I(N__3207));
    InMux I__509 (
            .O(N__3210),
            .I(N__3204));
    InMux I__508 (
            .O(N__3207),
            .I(N__3201));
    LocalMux I__507 (
            .O(N__3204),
            .I(N__3198));
    LocalMux I__506 (
            .O(N__3201),
            .I(\led_blink_inst.r_Count_2Z0Z_12 ));
    Odrv4 I__505 (
            .O(N__3198),
            .I(\led_blink_inst.r_Count_2Z0Z_12 ));
    InMux I__504 (
            .O(N__3193),
            .I(N__3190));
    LocalMux I__503 (
            .O(N__3190),
            .I(N__3187));
    Span4Mux_v I__502 (
            .O(N__3187),
            .I(N__3184));
    Odrv4 I__501 (
            .O(N__3184),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_12 ));
    InMux I__500 (
            .O(N__3181),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_11 ));
    InMux I__499 (
            .O(N__3178),
            .I(N__3175));
    LocalMux I__498 (
            .O(N__3175),
            .I(\led_blink_inst.o_LED_23_13 ));
    CascadeMux I__497 (
            .O(N__3172),
            .I(\led_blink_inst.o_LED_23_12_cascade_ ));
    InMux I__496 (
            .O(N__3169),
            .I(N__3166));
    LocalMux I__495 (
            .O(N__3166),
            .I(\led_blink_inst.o_LED_23_15 ));
    CascadeMux I__494 (
            .O(N__3163),
            .I(\led_blink_inst.o_LED_23_21_cascade_ ));
    InMux I__493 (
            .O(N__3160),
            .I(N__3154));
    InMux I__492 (
            .O(N__3159),
            .I(N__3154));
    LocalMux I__491 (
            .O(N__3154),
            .I(N__3150));
    InMux I__490 (
            .O(N__3153),
            .I(N__3147));
    Odrv4 I__489 (
            .O(N__3150),
            .I(\led_blink_inst.r_Count_2Z0Z_1 ));
    LocalMux I__488 (
            .O(N__3147),
            .I(\led_blink_inst.r_Count_2Z0Z_1 ));
    CascadeMux I__487 (
            .O(N__3142),
            .I(N__3138));
    CascadeMux I__486 (
            .O(N__3141),
            .I(N__3133));
    InMux I__485 (
            .O(N__3138),
            .I(N__3126));
    InMux I__484 (
            .O(N__3137),
            .I(N__3126));
    InMux I__483 (
            .O(N__3136),
            .I(N__3126));
    InMux I__482 (
            .O(N__3133),
            .I(N__3123));
    LocalMux I__481 (
            .O(N__3126),
            .I(\led_blink_inst.r_Count_2Z0Z_0 ));
    LocalMux I__480 (
            .O(N__3123),
            .I(\led_blink_inst.r_Count_2Z0Z_0 ));
    CascadeMux I__479 (
            .O(N__3118),
            .I(N__3114));
    CascadeMux I__478 (
            .O(N__3117),
            .I(N__3111));
    InMux I__477 (
            .O(N__3114),
            .I(N__3108));
    InMux I__476 (
            .O(N__3111),
            .I(N__3105));
    LocalMux I__475 (
            .O(N__3108),
            .I(\led_blink_inst.r_Count_2Z0Z_2 ));
    LocalMux I__474 (
            .O(N__3105),
            .I(\led_blink_inst.r_Count_2Z0Z_2 ));
    InMux I__473 (
            .O(N__3100),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_1 ));
    InMux I__472 (
            .O(N__3097),
            .I(N__3093));
    InMux I__471 (
            .O(N__3096),
            .I(N__3090));
    LocalMux I__470 (
            .O(N__3093),
            .I(\led_blink_inst.r_Count_2Z0Z_3 ));
    LocalMux I__469 (
            .O(N__3090),
            .I(\led_blink_inst.r_Count_2Z0Z_3 ));
    InMux I__468 (
            .O(N__3085),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_2 ));
    InMux I__467 (
            .O(N__3082),
            .I(N__3078));
    InMux I__466 (
            .O(N__3081),
            .I(N__3075));
    LocalMux I__465 (
            .O(N__3078),
            .I(\led_blink_inst.r_Count_2Z0Z_4 ));
    LocalMux I__464 (
            .O(N__3075),
            .I(\led_blink_inst.r_Count_2Z0Z_4 ));
    InMux I__463 (
            .O(N__3070),
            .I(N__3067));
    LocalMux I__462 (
            .O(N__3067),
            .I(\led_blink_inst.r_Count_2_RNO_0Z0Z_4 ));
    InMux I__461 (
            .O(N__3064),
            .I(\led_blink_inst.un2_r_Count_2_1_cry_3 ));
    CascadeMux I__460 (
            .O(N__3061),
            .I(N__3058));
    InMux I__459 (
            .O(N__3058),
            .I(N__3054));
    CascadeMux I__458 (
            .O(N__3057),
            .I(N__3051));
    LocalMux I__457 (
            .O(N__3054),
            .I(N__3048));
    InMux I__456 (
            .O(N__3051),
            .I(N__3045));
    Odrv4 I__455 (
            .O(N__3048),
            .I(\led_blink_inst.r_Count_1Z0Z_22 ));
    LocalMux I__454 (
            .O(N__3045),
            .I(\led_blink_inst.r_Count_1Z0Z_22 ));
    InMux I__453 (
            .O(N__3040),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_21 ));
    InMux I__452 (
            .O(N__3037),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_22 ));
    InMux I__451 (
            .O(N__3034),
            .I(N__3031));
    LocalMux I__450 (
            .O(N__3031),
            .I(N__3019));
    InMux I__449 (
            .O(N__3030),
            .I(N__3010));
    InMux I__448 (
            .O(N__3029),
            .I(N__3010));
    InMux I__447 (
            .O(N__3028),
            .I(N__3010));
    InMux I__446 (
            .O(N__3027),
            .I(N__3010));
    InMux I__445 (
            .O(N__3026),
            .I(N__2999));
    InMux I__444 (
            .O(N__3025),
            .I(N__2999));
    InMux I__443 (
            .O(N__3024),
            .I(N__2999));
    InMux I__442 (
            .O(N__3023),
            .I(N__2999));
    InMux I__441 (
            .O(N__3022),
            .I(N__2999));
    Span4Mux_v I__440 (
            .O(N__3019),
            .I(N__2992));
    LocalMux I__439 (
            .O(N__3010),
            .I(N__2989));
    LocalMux I__438 (
            .O(N__2999),
            .I(N__2986));
    InMux I__437 (
            .O(N__2998),
            .I(N__2977));
    InMux I__436 (
            .O(N__2997),
            .I(N__2977));
    InMux I__435 (
            .O(N__2996),
            .I(N__2977));
    InMux I__434 (
            .O(N__2995),
            .I(N__2977));
    Odrv4 I__433 (
            .O(N__2992),
            .I(\led_blink_inst.o_LED_13_17 ));
    Odrv12 I__432 (
            .O(N__2989),
            .I(\led_blink_inst.o_LED_13_17 ));
    Odrv4 I__431 (
            .O(N__2986),
            .I(\led_blink_inst.o_LED_13_17 ));
    LocalMux I__430 (
            .O(N__2977),
            .I(\led_blink_inst.o_LED_13_17 ));
    InMux I__429 (
            .O(N__2968),
            .I(N__2953));
    InMux I__428 (
            .O(N__2967),
            .I(N__2944));
    InMux I__427 (
            .O(N__2966),
            .I(N__2944));
    InMux I__426 (
            .O(N__2965),
            .I(N__2944));
    InMux I__425 (
            .O(N__2964),
            .I(N__2944));
    InMux I__424 (
            .O(N__2963),
            .I(N__2935));
    InMux I__423 (
            .O(N__2962),
            .I(N__2935));
    InMux I__422 (
            .O(N__2961),
            .I(N__2935));
    InMux I__421 (
            .O(N__2960),
            .I(N__2935));
    InMux I__420 (
            .O(N__2959),
            .I(N__2926));
    InMux I__419 (
            .O(N__2958),
            .I(N__2926));
    InMux I__418 (
            .O(N__2957),
            .I(N__2926));
    InMux I__417 (
            .O(N__2956),
            .I(N__2926));
    LocalMux I__416 (
            .O(N__2953),
            .I(\led_blink_inst.o_LED_13_16 ));
    LocalMux I__415 (
            .O(N__2944),
            .I(\led_blink_inst.o_LED_13_16 ));
    LocalMux I__414 (
            .O(N__2935),
            .I(\led_blink_inst.o_LED_13_16 ));
    LocalMux I__413 (
            .O(N__2926),
            .I(\led_blink_inst.o_LED_13_16 ));
    CascadeMux I__412 (
            .O(N__2917),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_23_cascade_ ));
    CascadeMux I__411 (
            .O(N__2914),
            .I(N__2903));
    CascadeMux I__410 (
            .O(N__2913),
            .I(N__2900));
    CascadeMux I__409 (
            .O(N__2912),
            .I(N__2897));
    CascadeMux I__408 (
            .O(N__2911),
            .I(N__2892));
    CascadeMux I__407 (
            .O(N__2910),
            .I(N__2887));
    CascadeMux I__406 (
            .O(N__2909),
            .I(N__2884));
    CascadeMux I__405 (
            .O(N__2908),
            .I(N__2881));
    InMux I__404 (
            .O(N__2907),
            .I(N__2878));
    InMux I__403 (
            .O(N__2906),
            .I(N__2869));
    InMux I__402 (
            .O(N__2903),
            .I(N__2869));
    InMux I__401 (
            .O(N__2900),
            .I(N__2869));
    InMux I__400 (
            .O(N__2897),
            .I(N__2869));
    InMux I__399 (
            .O(N__2896),
            .I(N__2860));
    InMux I__398 (
            .O(N__2895),
            .I(N__2860));
    InMux I__397 (
            .O(N__2892),
            .I(N__2860));
    InMux I__396 (
            .O(N__2891),
            .I(N__2860));
    InMux I__395 (
            .O(N__2890),
            .I(N__2851));
    InMux I__394 (
            .O(N__2887),
            .I(N__2851));
    InMux I__393 (
            .O(N__2884),
            .I(N__2851));
    InMux I__392 (
            .O(N__2881),
            .I(N__2851));
    LocalMux I__391 (
            .O(N__2878),
            .I(\led_blink_inst.o_LED_13_21 ));
    LocalMux I__390 (
            .O(N__2869),
            .I(\led_blink_inst.o_LED_13_21 ));
    LocalMux I__389 (
            .O(N__2860),
            .I(\led_blink_inst.o_LED_13_21 ));
    LocalMux I__388 (
            .O(N__2851),
            .I(\led_blink_inst.o_LED_13_21 ));
    CascadeMux I__387 (
            .O(N__2842),
            .I(N__2839));
    InMux I__386 (
            .O(N__2839),
            .I(N__2836));
    LocalMux I__385 (
            .O(N__2836),
            .I(N__2832));
    InMux I__384 (
            .O(N__2835),
            .I(N__2829));
    Odrv4 I__383 (
            .O(N__2832),
            .I(\led_blink_inst.r_Count_1Z0Z_23 ));
    LocalMux I__382 (
            .O(N__2829),
            .I(\led_blink_inst.r_Count_1Z0Z_23 ));
    IoInMux I__381 (
            .O(N__2824),
            .I(N__2821));
    LocalMux I__380 (
            .O(N__2821),
            .I(N__2817));
    CascadeMux I__379 (
            .O(N__2820),
            .I(N__2814));
    Span4Mux_s3_h I__378 (
            .O(N__2817),
            .I(N__2811));
    InMux I__377 (
            .O(N__2814),
            .I(N__2808));
    Odrv4 I__376 (
            .O(N__2811),
            .I(o_LED_2_c));
    LocalMux I__375 (
            .O(N__2808),
            .I(o_LED_2_c));
    InMux I__374 (
            .O(N__2803),
            .I(N__2800));
    LocalMux I__373 (
            .O(N__2800),
            .I(N__2797));
    Odrv4 I__372 (
            .O(N__2797),
            .I(\led_blink_inst.o_LED_23_14 ));
    CascadeMux I__371 (
            .O(N__2794),
            .I(N__2790));
    CascadeMux I__370 (
            .O(N__2793),
            .I(N__2787));
    InMux I__369 (
            .O(N__2790),
            .I(N__2784));
    InMux I__368 (
            .O(N__2787),
            .I(N__2781));
    LocalMux I__367 (
            .O(N__2784),
            .I(\led_blink_inst.r_Count_1Z0Z_14 ));
    LocalMux I__366 (
            .O(N__2781),
            .I(\led_blink_inst.r_Count_1Z0Z_14 ));
    InMux I__365 (
            .O(N__2776),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_13 ));
    CascadeMux I__364 (
            .O(N__2773),
            .I(N__2769));
    InMux I__363 (
            .O(N__2772),
            .I(N__2766));
    InMux I__362 (
            .O(N__2769),
            .I(N__2763));
    LocalMux I__361 (
            .O(N__2766),
            .I(\led_blink_inst.r_Count_1Z0Z_15 ));
    LocalMux I__360 (
            .O(N__2763),
            .I(\led_blink_inst.r_Count_1Z0Z_15 ));
    CascadeMux I__359 (
            .O(N__2758),
            .I(N__2755));
    InMux I__358 (
            .O(N__2755),
            .I(N__2752));
    LocalMux I__357 (
            .O(N__2752),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_15 ));
    InMux I__356 (
            .O(N__2749),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_14 ));
    InMux I__355 (
            .O(N__2746),
            .I(N__2742));
    CascadeMux I__354 (
            .O(N__2745),
            .I(N__2739));
    LocalMux I__353 (
            .O(N__2742),
            .I(N__2736));
    InMux I__352 (
            .O(N__2739),
            .I(N__2733));
    Odrv4 I__351 (
            .O(N__2736),
            .I(\led_blink_inst.r_Count_1Z0Z_16 ));
    LocalMux I__350 (
            .O(N__2733),
            .I(\led_blink_inst.r_Count_1Z0Z_16 ));
    InMux I__349 (
            .O(N__2728),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_15 ));
    CascadeMux I__348 (
            .O(N__2725),
            .I(N__2721));
    InMux I__347 (
            .O(N__2724),
            .I(N__2718));
    InMux I__346 (
            .O(N__2721),
            .I(N__2715));
    LocalMux I__345 (
            .O(N__2718),
            .I(\led_blink_inst.r_Count_1Z0Z_17 ));
    LocalMux I__344 (
            .O(N__2715),
            .I(\led_blink_inst.r_Count_1Z0Z_17 ));
    InMux I__343 (
            .O(N__2710),
            .I(N__2707));
    LocalMux I__342 (
            .O(N__2707),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_17 ));
    InMux I__341 (
            .O(N__2704),
            .I(bfn_8_9_0_));
    CascadeMux I__340 (
            .O(N__2701),
            .I(N__2697));
    InMux I__339 (
            .O(N__2700),
            .I(N__2694));
    InMux I__338 (
            .O(N__2697),
            .I(N__2691));
    LocalMux I__337 (
            .O(N__2694),
            .I(\led_blink_inst.r_Count_1Z0Z_18 ));
    LocalMux I__336 (
            .O(N__2691),
            .I(\led_blink_inst.r_Count_1Z0Z_18 ));
    InMux I__335 (
            .O(N__2686),
            .I(N__2683));
    LocalMux I__334 (
            .O(N__2683),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_18 ));
    InMux I__333 (
            .O(N__2680),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_17 ));
    CascadeMux I__332 (
            .O(N__2677),
            .I(N__2673));
    InMux I__331 (
            .O(N__2676),
            .I(N__2670));
    InMux I__330 (
            .O(N__2673),
            .I(N__2667));
    LocalMux I__329 (
            .O(N__2670),
            .I(\led_blink_inst.r_Count_1Z0Z_19 ));
    LocalMux I__328 (
            .O(N__2667),
            .I(\led_blink_inst.r_Count_1Z0Z_19 ));
    InMux I__327 (
            .O(N__2662),
            .I(N__2659));
    LocalMux I__326 (
            .O(N__2659),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_19 ));
    InMux I__325 (
            .O(N__2656),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_18 ));
    CascadeMux I__324 (
            .O(N__2653),
            .I(N__2649));
    InMux I__323 (
            .O(N__2652),
            .I(N__2646));
    InMux I__322 (
            .O(N__2649),
            .I(N__2643));
    LocalMux I__321 (
            .O(N__2646),
            .I(\led_blink_inst.r_Count_1Z0Z_20 ));
    LocalMux I__320 (
            .O(N__2643),
            .I(\led_blink_inst.r_Count_1Z0Z_20 ));
    InMux I__319 (
            .O(N__2638),
            .I(N__2635));
    LocalMux I__318 (
            .O(N__2635),
            .I(N__2632));
    Span4Mux_h I__317 (
            .O(N__2632),
            .I(N__2629));
    Odrv4 I__316 (
            .O(N__2629),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_20 ));
    InMux I__315 (
            .O(N__2626),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_19 ));
    CascadeMux I__314 (
            .O(N__2623),
            .I(N__2619));
    InMux I__313 (
            .O(N__2622),
            .I(N__2616));
    InMux I__312 (
            .O(N__2619),
            .I(N__2613));
    LocalMux I__311 (
            .O(N__2616),
            .I(\led_blink_inst.r_Count_1Z0Z_21 ));
    LocalMux I__310 (
            .O(N__2613),
            .I(\led_blink_inst.r_Count_1Z0Z_21 ));
    CascadeMux I__309 (
            .O(N__2608),
            .I(N__2605));
    InMux I__308 (
            .O(N__2605),
            .I(N__2602));
    LocalMux I__307 (
            .O(N__2602),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_21 ));
    InMux I__306 (
            .O(N__2599),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_20 ));
    InMux I__305 (
            .O(N__2596),
            .I(N__2592));
    InMux I__304 (
            .O(N__2595),
            .I(N__2589));
    LocalMux I__303 (
            .O(N__2592),
            .I(\led_blink_inst.r_Count_1Z0Z_6 ));
    LocalMux I__302 (
            .O(N__2589),
            .I(\led_blink_inst.r_Count_1Z0Z_6 ));
    InMux I__301 (
            .O(N__2584),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_5 ));
    InMux I__300 (
            .O(N__2581),
            .I(N__2578));
    LocalMux I__299 (
            .O(N__2578),
            .I(N__2575));
    Span4Mux_v I__298 (
            .O(N__2575),
            .I(N__2571));
    InMux I__297 (
            .O(N__2574),
            .I(N__2568));
    Odrv4 I__296 (
            .O(N__2571),
            .I(\led_blink_inst.r_Count_1Z0Z_7 ));
    LocalMux I__295 (
            .O(N__2568),
            .I(\led_blink_inst.r_Count_1Z0Z_7 ));
    InMux I__294 (
            .O(N__2563),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_6 ));
    CascadeMux I__293 (
            .O(N__2560),
            .I(N__2556));
    InMux I__292 (
            .O(N__2559),
            .I(N__2553));
    InMux I__291 (
            .O(N__2556),
            .I(N__2550));
    LocalMux I__290 (
            .O(N__2553),
            .I(\led_blink_inst.r_Count_1Z0Z_8 ));
    LocalMux I__289 (
            .O(N__2550),
            .I(\led_blink_inst.r_Count_1Z0Z_8 ));
    InMux I__288 (
            .O(N__2545),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_7 ));
    CascadeMux I__287 (
            .O(N__2542),
            .I(N__2538));
    InMux I__286 (
            .O(N__2541),
            .I(N__2535));
    InMux I__285 (
            .O(N__2538),
            .I(N__2532));
    LocalMux I__284 (
            .O(N__2535),
            .I(\led_blink_inst.r_Count_1Z0Z_9 ));
    LocalMux I__283 (
            .O(N__2532),
            .I(\led_blink_inst.r_Count_1Z0Z_9 ));
    InMux I__282 (
            .O(N__2527),
            .I(bfn_8_8_0_));
    InMux I__281 (
            .O(N__2524),
            .I(N__2520));
    InMux I__280 (
            .O(N__2523),
            .I(N__2517));
    LocalMux I__279 (
            .O(N__2520),
            .I(\led_blink_inst.r_Count_1Z0Z_10 ));
    LocalMux I__278 (
            .O(N__2517),
            .I(\led_blink_inst.r_Count_1Z0Z_10 ));
    CascadeMux I__277 (
            .O(N__2512),
            .I(N__2509));
    InMux I__276 (
            .O(N__2509),
            .I(N__2506));
    LocalMux I__275 (
            .O(N__2506),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_10 ));
    InMux I__274 (
            .O(N__2503),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_9 ));
    CascadeMux I__273 (
            .O(N__2500),
            .I(N__2497));
    InMux I__272 (
            .O(N__2497),
            .I(N__2493));
    InMux I__271 (
            .O(N__2496),
            .I(N__2490));
    LocalMux I__270 (
            .O(N__2493),
            .I(\led_blink_inst.r_Count_1Z0Z_11 ));
    LocalMux I__269 (
            .O(N__2490),
            .I(\led_blink_inst.r_Count_1Z0Z_11 ));
    InMux I__268 (
            .O(N__2485),
            .I(N__2482));
    LocalMux I__267 (
            .O(N__2482),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_11 ));
    InMux I__266 (
            .O(N__2479),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_10 ));
    CascadeMux I__265 (
            .O(N__2476),
            .I(N__2472));
    InMux I__264 (
            .O(N__2475),
            .I(N__2469));
    InMux I__263 (
            .O(N__2472),
            .I(N__2466));
    LocalMux I__262 (
            .O(N__2469),
            .I(\led_blink_inst.r_Count_1Z0Z_12 ));
    LocalMux I__261 (
            .O(N__2466),
            .I(\led_blink_inst.r_Count_1Z0Z_12 ));
    InMux I__260 (
            .O(N__2461),
            .I(N__2458));
    LocalMux I__259 (
            .O(N__2458),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_12 ));
    InMux I__258 (
            .O(N__2455),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_11 ));
    CascadeMux I__257 (
            .O(N__2452),
            .I(N__2448));
    InMux I__256 (
            .O(N__2451),
            .I(N__2445));
    InMux I__255 (
            .O(N__2448),
            .I(N__2442));
    LocalMux I__254 (
            .O(N__2445),
            .I(\led_blink_inst.r_Count_1Z0Z_13 ));
    LocalMux I__253 (
            .O(N__2442),
            .I(\led_blink_inst.r_Count_1Z0Z_13 ));
    CascadeMux I__252 (
            .O(N__2437),
            .I(N__2434));
    InMux I__251 (
            .O(N__2434),
            .I(N__2431));
    LocalMux I__250 (
            .O(N__2431),
            .I(N__2428));
    Odrv4 I__249 (
            .O(N__2428),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_13 ));
    InMux I__248 (
            .O(N__2425),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_12 ));
    InMux I__247 (
            .O(N__2422),
            .I(N__2417));
    InMux I__246 (
            .O(N__2421),
            .I(N__2414));
    InMux I__245 (
            .O(N__2420),
            .I(N__2411));
    LocalMux I__244 (
            .O(N__2417),
            .I(\led_blink_inst.r_Count_1Z0Z_1 ));
    LocalMux I__243 (
            .O(N__2414),
            .I(\led_blink_inst.r_Count_1Z0Z_1 ));
    LocalMux I__242 (
            .O(N__2411),
            .I(\led_blink_inst.r_Count_1Z0Z_1 ));
    CascadeMux I__241 (
            .O(N__2404),
            .I(N__2398));
    InMux I__240 (
            .O(N__2403),
            .I(N__2395));
    InMux I__239 (
            .O(N__2402),
            .I(N__2392));
    InMux I__238 (
            .O(N__2401),
            .I(N__2389));
    InMux I__237 (
            .O(N__2398),
            .I(N__2386));
    LocalMux I__236 (
            .O(N__2395),
            .I(\led_blink_inst.r_Count_1Z0Z_0 ));
    LocalMux I__235 (
            .O(N__2392),
            .I(\led_blink_inst.r_Count_1Z0Z_0 ));
    LocalMux I__234 (
            .O(N__2389),
            .I(\led_blink_inst.r_Count_1Z0Z_0 ));
    LocalMux I__233 (
            .O(N__2386),
            .I(\led_blink_inst.r_Count_1Z0Z_0 ));
    CascadeMux I__232 (
            .O(N__2377),
            .I(N__2374));
    InMux I__231 (
            .O(N__2374),
            .I(N__2370));
    InMux I__230 (
            .O(N__2373),
            .I(N__2367));
    LocalMux I__229 (
            .O(N__2370),
            .I(\led_blink_inst.r_Count_1Z0Z_2 ));
    LocalMux I__228 (
            .O(N__2367),
            .I(\led_blink_inst.r_Count_1Z0Z_2 ));
    InMux I__227 (
            .O(N__2362),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_1 ));
    InMux I__226 (
            .O(N__2359),
            .I(N__2355));
    InMux I__225 (
            .O(N__2358),
            .I(N__2352));
    LocalMux I__224 (
            .O(N__2355),
            .I(\led_blink_inst.r_Count_1Z0Z_3 ));
    LocalMux I__223 (
            .O(N__2352),
            .I(\led_blink_inst.r_Count_1Z0Z_3 ));
    InMux I__222 (
            .O(N__2347),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_2 ));
    CascadeMux I__221 (
            .O(N__2344),
            .I(N__2340));
    InMux I__220 (
            .O(N__2343),
            .I(N__2337));
    InMux I__219 (
            .O(N__2340),
            .I(N__2334));
    LocalMux I__218 (
            .O(N__2337),
            .I(\led_blink_inst.r_Count_1Z0Z_4 ));
    LocalMux I__217 (
            .O(N__2334),
            .I(\led_blink_inst.r_Count_1Z0Z_4 ));
    InMux I__216 (
            .O(N__2329),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_3 ));
    InMux I__215 (
            .O(N__2326),
            .I(N__2322));
    InMux I__214 (
            .O(N__2325),
            .I(N__2319));
    LocalMux I__213 (
            .O(N__2322),
            .I(\led_blink_inst.r_Count_1Z0Z_5 ));
    LocalMux I__212 (
            .O(N__2319),
            .I(\led_blink_inst.r_Count_1Z0Z_5 ));
    InMux I__211 (
            .O(N__2314),
            .I(N__2311));
    LocalMux I__210 (
            .O(N__2311),
            .I(\led_blink_inst.r_Count_1_RNO_0Z0Z_5 ));
    InMux I__209 (
            .O(N__2308),
            .I(\led_blink_inst.un3_r_Count_1_1_cry_4 ));
    CascadeMux I__208 (
            .O(N__2305),
            .I(\led_blink_inst.o_LED_23_16_cascade_ ));
    InMux I__207 (
            .O(N__2302),
            .I(N__2299));
    LocalMux I__206 (
            .O(N__2299),
            .I(\led_blink_inst.o_LED_13_15 ));
    InMux I__205 (
            .O(N__2296),
            .I(N__2293));
    LocalMux I__204 (
            .O(N__2293),
            .I(\led_blink_inst.o_LED_13_13 ));
    CascadeMux I__203 (
            .O(N__2290),
            .I(\led_blink_inst.o_LED_13_14_cascade_ ));
    InMux I__202 (
            .O(N__2287),
            .I(N__2284));
    LocalMux I__201 (
            .O(N__2284),
            .I(\led_blink_inst.o_LED_13_12 ));
    CascadeMux I__200 (
            .O(N__2281),
            .I(\led_blink_inst.o_LED_13_21_cascade_ ));
    CascadeMux I__199 (
            .O(N__2278),
            .I(\led_blink_inst.o_LED_13_16_cascade_ ));
    IoInMux I__198 (
            .O(N__2275),
            .I(N__2272));
    LocalMux I__197 (
            .O(N__2272),
            .I(N__2269));
    IoSpan4Mux I__196 (
            .O(N__2269),
            .I(N__2266));
    Span4Mux_s3_h I__195 (
            .O(N__2266),
            .I(N__2262));
    InMux I__194 (
            .O(N__2265),
            .I(N__2259));
    Odrv4 I__193 (
            .O(N__2262),
            .I(o_LED_1_c));
    LocalMux I__192 (
            .O(N__2259),
            .I(o_LED_1_c));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\led_blink_inst.un3_r_Count_1_1_cry_8 ),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\led_blink_inst.un3_r_Count_1_1_cry_16 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(\led_blink_inst.un2_r_Count_4_1_cry_8 ),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\led_blink_inst.un2_r_Count_4_1_cry_16 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_12_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_3_0_));
    defparam IN_MUX_bfv_12_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_4_0_ (
            .carryinitin(\led_blink_inst.un2_r_Count_3_1_cry_8 ),
            .carryinitout(bfn_12_4_0_));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(\led_blink_inst.un2_r_Count_3_1_cry_16 ),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(\led_blink_inst.un2_r_Count_2_1_cry_8 ),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(\led_blink_inst.un2_r_Count_2_1_cry_16 ),
            .carryinitout(bfn_9_8_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNIVTTA_13_LC_6_8_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_RNIVTTA_13_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNIVTTA_13_LC_6_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_1_RNIVTTA_13_LC_6_8_7  (
            .in0(N__2772),
            .in1(N__2451),
            .in2(N__2701),
            .in3(N__2724),
            .lcout(\led_blink_inst.o_LED_13_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNIJ5RV_16_LC_7_6_0 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_RNIJ5RV_16_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNIJ5RV_16_LC_7_6_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_1_RNIJ5RV_16_LC_7_6_0  (
            .in0(N__2746),
            .in1(N__2343),
            .in2(N__3061),
            .in3(N__2401),
            .lcout(\led_blink_inst.o_LED_13_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_0_LC_7_7_0 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_0_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_0_LC_7_7_0 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \led_blink_inst.r_Count_1_0_LC_7_7_0  (
            .in0(N__2996),
            .in1(N__2957),
            .in2(N__2909),
            .in3(N__2402),
            .lcout(\led_blink_inst.r_Count_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4929),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNILPMK1_1_LC_7_7_1 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_RNILPMK1_1_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNILPMK1_1_LC_7_7_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_1_RNILPMK1_1_LC_7_7_1  (
            .in0(N__2421),
            .in1(N__2596),
            .in2(N__2377),
            .in3(N__2559),
            .lcout(\led_blink_inst.o_LED_13_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNICN8A1_14_LC_7_7_3 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_RNICN8A1_14_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNICN8A1_14_LC_7_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_1_RNICN8A1_14_LC_7_7_3  (
            .in0(N__2581),
            .in1(N__2359),
            .in2(N__2794),
            .in3(N__2541),
            .lcout(\led_blink_inst.o_LED_13_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.o_LED_1_LC_7_7_4 .C_ON=1'b0;
    defparam \led_blink_inst.o_LED_1_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.o_LED_1_LC_7_7_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \led_blink_inst.o_LED_1_LC_7_7_4  (
            .in0(N__2995),
            .in1(N__2265),
            .in2(N__2908),
            .in3(N__2956),
            .lcout(o_LED_1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4929),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_5_LC_7_7_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_5_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_5_LC_7_7_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_1_5_LC_7_7_6  (
            .in0(N__2998),
            .in1(N__2959),
            .in2(N__2910),
            .in3(N__2314),
            .lcout(\led_blink_inst.r_Count_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4929),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_15_LC_7_7_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_15_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_15_LC_7_7_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_1_15_LC_7_7_7  (
            .in0(N__2958),
            .in1(N__2997),
            .in2(N__2758),
            .in3(N__2890),
            .lcout(\led_blink_inst.r_Count_1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4929),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNIVMBL_10_LC_7_8_0 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_RNIVMBL_10_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNIVMBL_10_LC_7_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_1_RNIVMBL_10_LC_7_8_0  (
            .in0(N__2524),
            .in1(N__2326),
            .in2(N__2500),
            .in3(N__2475),
            .lcout(),
            .ltout(\led_blink_inst.o_LED_13_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNIV59V3_10_LC_7_8_1 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_RNIV59V3_10_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNIV59V3_10_LC_7_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_1_RNIV59V3_10_LC_7_8_1  (
            .in0(N__2302),
            .in1(N__2296),
            .in2(N__2290),
            .in3(N__2287),
            .lcout(\led_blink_inst.o_LED_13_21 ),
            .ltout(\led_blink_inst.o_LED_13_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_20_LC_7_8_2 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_20_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_20_LC_7_8_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_1_20_LC_7_8_2  (
            .in0(N__2963),
            .in1(N__3026),
            .in2(N__2281),
            .in3(N__2638),
            .lcout(\led_blink_inst.r_Count_1Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4927),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNIOP0B_23_LC_7_8_3 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_RNIOP0B_23_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNIOP0B_23_LC_7_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_1_RNIOP0B_23_LC_7_8_3  (
            .in0(N__2622),
            .in1(N__2652),
            .in2(N__2842),
            .in3(N__2676),
            .lcout(\led_blink_inst.o_LED_13_16 ),
            .ltout(\led_blink_inst.o_LED_13_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_11_LC_7_8_4 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_11_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_11_LC_7_8_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_1_11_LC_7_8_4  (
            .in0(N__2891),
            .in1(N__3023),
            .in2(N__2278),
            .in3(N__2485),
            .lcout(\led_blink_inst.r_Count_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4927),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_13_LC_7_8_5 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_13_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_13_LC_7_8_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_1_13_LC_7_8_5  (
            .in0(N__3025),
            .in1(N__2962),
            .in2(N__2437),
            .in3(N__2896),
            .lcout(\led_blink_inst.r_Count_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4927),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_12_LC_7_8_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_12_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_12_LC_7_8_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_1_12_LC_7_8_6  (
            .in0(N__2961),
            .in1(N__3024),
            .in2(N__2911),
            .in3(N__2461),
            .lcout(\led_blink_inst.r_Count_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4927),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_10_LC_7_8_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_10_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_10_LC_7_8_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_1_10_LC_7_8_7  (
            .in0(N__3022),
            .in1(N__2960),
            .in2(N__2512),
            .in3(N__2895),
            .lcout(\led_blink_inst.r_Count_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4927),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_18_LC_7_9_0 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_18_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_18_LC_7_9_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_1_18_LC_7_9_0  (
            .in0(N__3028),
            .in1(N__2965),
            .in2(N__2913),
            .in3(N__2686),
            .lcout(\led_blink_inst.r_Count_1Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4930),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_17_LC_7_9_2 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_17_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_17_LC_7_9_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_1_17_LC_7_9_2  (
            .in0(N__3027),
            .in1(N__2964),
            .in2(N__2912),
            .in3(N__2710),
            .lcout(\led_blink_inst.r_Count_1Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4930),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_19_LC_7_9_4 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_19_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_19_LC_7_9_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_1_19_LC_7_9_4  (
            .in0(N__3029),
            .in1(N__2966),
            .in2(N__2914),
            .in3(N__2662),
            .lcout(\led_blink_inst.r_Count_1Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4930),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_21_LC_7_9_5 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_21_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_21_LC_7_9_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_1_21_LC_7_9_5  (
            .in0(N__2967),
            .in1(N__3030),
            .in2(N__2608),
            .in3(N__2906),
            .lcout(\led_blink_inst.r_Count_1Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4930),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNI1EOR_18_LC_8_5_1 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_RNI1EOR_18_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNI1EOR_18_LC_8_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_2_RNI1EOR_18_LC_8_5_1  (
            .in0(N__3393),
            .in1(N__3426),
            .in2(N__3604),
            .in3(N__3453),
            .lcout(\led_blink_inst.o_LED_23_16 ),
            .ltout(\led_blink_inst.o_LED_23_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_12_LC_8_5_2 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_12_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_12_LC_8_5_2 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \led_blink_inst.r_Count_2_12_LC_8_5_2  (
            .in0(N__3193),
            .in1(N__3791),
            .in2(N__2305),
            .in3(N__3655),
            .lcout(\led_blink_inst.r_Count_2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4937),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNIOJCA1_10_LC_8_5_5 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_RNIOJCA1_10_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNIOJCA1_10_LC_8_5_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_2_RNIOJCA1_10_LC_8_5_5  (
            .in0(N__3301),
            .in1(N__3082),
            .in2(N__3244),
            .in3(N__3270),
            .lcout(\led_blink_inst.o_LED_23_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNIV9MR_12_LC_8_5_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_RNIV9MR_12_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNIV9MR_12_LC_8_5_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_2_RNIV9MR_12_LC_8_5_6  (
            .in0(N__3562),
            .in1(N__3519),
            .in2(N__3211),
            .in3(N__3489),
            .lcout(\led_blink_inst.o_LED_23_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_17_LC_8_6_0 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_17_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_17_LC_8_6_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_2_17_LC_8_6_0  (
            .in0(N__3794),
            .in1(N__3729),
            .in2(N__3475),
            .in3(N__3660),
            .lcout(\led_blink_inst.r_Count_2Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4934),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_1_LC_8_6_1 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_1_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_1_LC_8_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \led_blink_inst.r_Count_1_1_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__2403),
            .in2(_gnd_net_),
            .in3(N__2422),
            .lcout(\led_blink_inst.r_Count_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4934),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_20_LC_8_6_2 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_20_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_20_LC_8_6_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_2_20_LC_8_6_2  (
            .in0(N__3797),
            .in1(N__3732),
            .in2(N__3379),
            .in3(N__3665),
            .lcout(\led_blink_inst.r_Count_2Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4934),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_19_LC_8_6_4 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_19_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_19_LC_8_6_4 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_2_19_LC_8_6_4  (
            .in0(N__3796),
            .in1(N__3731),
            .in2(N__3412),
            .in3(N__3664),
            .lcout(\led_blink_inst.r_Count_2Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4934),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_18_LC_8_6_5 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_18_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_18_LC_8_6_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_2_18_LC_8_6_5  (
            .in0(N__3730),
            .in1(N__3795),
            .in2(N__3672),
            .in3(N__3439),
            .lcout(\led_blink_inst.r_Count_2Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4934),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_10_LC_8_6_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_10_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_10_LC_8_6_6 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_2_10_LC_8_6_6  (
            .in0(N__3792),
            .in1(N__3727),
            .in2(N__3256),
            .in3(N__3656),
            .lcout(\led_blink_inst.r_Count_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4934),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_14_LC_8_6_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_14_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_14_LC_8_6_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_2_14_LC_8_6_7  (
            .in0(N__3728),
            .in1(N__3793),
            .in2(N__3671),
            .in3(N__3550),
            .lcout(\led_blink_inst.r_Count_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4934),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.un3_r_Count_1_1_cry_1_c_LC_8_7_0 .C_ON=1'b1;
    defparam \led_blink_inst.un3_r_Count_1_1_cry_1_c_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.un3_r_Count_1_1_cry_1_c_LC_8_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \led_blink_inst.un3_r_Count_1_1_cry_1_c_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__2420),
            .in2(N__2404),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_2_LC_8_7_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_2_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_2_LC_8_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_1_2_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__2373),
            .in2(_gnd_net_),
            .in3(N__2362),
            .lcout(\led_blink_inst.r_Count_1Z0Z_2 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_1 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_2 ),
            .clk(N__4932),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_3_LC_8_7_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_3_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_3_LC_8_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_1_3_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__2358),
            .in2(_gnd_net_),
            .in3(N__2347),
            .lcout(\led_blink_inst.r_Count_1Z0Z_3 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_2 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_3 ),
            .clk(N__4932),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_4_LC_8_7_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_4_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_4_LC_8_7_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_4_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2344),
            .in3(N__2329),
            .lcout(\led_blink_inst.r_Count_1Z0Z_4 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_3 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_4 ),
            .clk(N__4932),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_5_LC_8_7_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_RNO_0_5_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_5_LC_8_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_5_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__2325),
            .in2(_gnd_net_),
            .in3(N__2308),
            .lcout(\led_blink_inst.r_Count_1_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_4 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_6_LC_8_7_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_6_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_6_LC_8_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_1_6_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__2595),
            .in2(_gnd_net_),
            .in3(N__2584),
            .lcout(\led_blink_inst.r_Count_1Z0Z_6 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_5 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_6 ),
            .clk(N__4932),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_7_LC_8_7_6 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_7_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_7_LC_8_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_1_7_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__2574),
            .in2(_gnd_net_),
            .in3(N__2563),
            .lcout(\led_blink_inst.r_Count_1Z0Z_7 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_6 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_7 ),
            .clk(N__4932),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_8_LC_8_7_7 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_8_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_8_LC_8_7_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_8_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2560),
            .in3(N__2545),
            .lcout(\led_blink_inst.r_Count_1Z0Z_8 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_7 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_8 ),
            .clk(N__4932),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_9_LC_8_8_0 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_9_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_9_LC_8_8_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_9_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2542),
            .in3(N__2527),
            .lcout(\led_blink_inst.r_Count_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_9 ),
            .clk(N__4928),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_10_LC_8_8_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_RNO_0_10_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_10_LC_8_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_10_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__2523),
            .in2(_gnd_net_),
            .in3(N__2503),
            .lcout(\led_blink_inst.r_Count_1_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_9 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_11_LC_8_8_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_RNO_0_11_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_11_LC_8_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_11_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__2496),
            .in2(_gnd_net_),
            .in3(N__2479),
            .lcout(\led_blink_inst.r_Count_1_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_10 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_12_LC_8_8_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_RNO_0_12_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_12_LC_8_8_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_12_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2476),
            .in3(N__2455),
            .lcout(\led_blink_inst.r_Count_1_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_11 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_13_LC_8_8_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_RNO_0_13_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_13_LC_8_8_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_13_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2452),
            .in3(N__2425),
            .lcout(\led_blink_inst.r_Count_1_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_12 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_14_LC_8_8_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_14_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_14_LC_8_8_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_14_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2793),
            .in3(N__2776),
            .lcout(\led_blink_inst.r_Count_1Z0Z_14 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_13 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_14 ),
            .clk(N__4928),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_15_LC_8_8_6 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_RNO_0_15_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_15_LC_8_8_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_15_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2773),
            .in3(N__2749),
            .lcout(\led_blink_inst.r_Count_1_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_14 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_16_LC_8_8_7 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_16_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_16_LC_8_8_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_16_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2745),
            .in3(N__2728),
            .lcout(\led_blink_inst.r_Count_1Z0Z_16 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_15 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_16 ),
            .clk(N__4928),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_17_LC_8_9_0 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_RNO_0_17_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_17_LC_8_9_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_17_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2725),
            .in3(N__2704),
            .lcout(\led_blink_inst.r_Count_1_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_18_LC_8_9_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_RNO_0_18_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_18_LC_8_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_18_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__2700),
            .in2(_gnd_net_),
            .in3(N__2680),
            .lcout(\led_blink_inst.r_Count_1_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_17 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_19_LC_8_9_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_RNO_0_19_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_19_LC_8_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_19_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2677),
            .in3(N__2656),
            .lcout(\led_blink_inst.r_Count_1_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_18 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_20_LC_8_9_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_RNO_0_20_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_20_LC_8_9_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_20_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2653),
            .in3(N__2626),
            .lcout(\led_blink_inst.r_Count_1_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_19 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_21_LC_8_9_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_RNO_0_21_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_21_LC_8_9_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_21_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2623),
            .in3(N__2599),
            .lcout(\led_blink_inst.r_Count_1_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_20 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_22_LC_8_9_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_1_22_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_22_LC_8_9_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_1_22_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3057),
            .in3(N__3040),
            .lcout(\led_blink_inst.r_Count_1Z0Z_22 ),
            .ltout(),
            .carryin(\led_blink_inst.un3_r_Count_1_1_cry_21 ),
            .carryout(\led_blink_inst.un3_r_Count_1_1_cry_22 ),
            .clk(N__4933),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_RNO_0_23_LC_8_9_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_RNO_0_23_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_1_RNO_0_23_LC_8_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \led_blink_inst.r_Count_1_RNO_0_23_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__2835),
            .in2(_gnd_net_),
            .in3(N__3037),
            .lcout(),
            .ltout(\led_blink_inst.r_Count_1_RNO_0Z0Z_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_1_23_LC_8_9_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_1_23_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_1_23_LC_8_9_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_1_23_LC_8_9_7  (
            .in0(N__3034),
            .in1(N__2968),
            .in2(N__2917),
            .in3(N__2907),
            .lcout(\led_blink_inst.r_Count_1Z0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4933),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_11_LC_9_4_3 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_11_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_11_LC_9_4_3 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_2_11_LC_9_4_3  (
            .in0(N__3725),
            .in1(N__3789),
            .in2(N__3226),
            .in3(N__3651),
            .lcout(\led_blink_inst.r_Count_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4944),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_16_LC_9_4_4 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_16_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_16_LC_9_4_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_2_16_LC_9_4_4  (
            .in0(N__3790),
            .in1(N__3726),
            .in2(N__3670),
            .in3(N__3505),
            .lcout(\led_blink_inst.r_Count_2Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4944),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.o_LED_2_LC_9_4_7 .C_ON=1'b0;
    defparam \led_blink_inst.o_LED_2_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.o_LED_2_LC_9_4_7 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \led_blink_inst.o_LED_2_LC_9_4_7  (
            .in0(N__3724),
            .in1(N__3788),
            .in2(N__2820),
            .in3(N__3650),
            .lcout(o_LED_2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4944),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_1_LC_9_5_0 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_1_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_1_LC_9_5_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_2_1_LC_9_5_0  (
            .in0(N__3160),
            .in1(_gnd_net_),
            .in2(N__3142),
            .in3(_gnd_net_),
            .lcout(\led_blink_inst.r_Count_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4941),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNI0SCA1_13_LC_9_5_1 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_RNI0SCA1_13_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNI0SCA1_13_LC_9_5_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_2_RNI0SCA1_13_LC_9_5_1  (
            .in0(N__3349),
            .in1(N__3316),
            .in2(N__3583),
            .in3(N__3541),
            .lcout(\led_blink_inst.o_LED_23_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNI7SOH1_23_LC_9_5_2 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_RNI7SOH1_23_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNI7SOH1_23_LC_9_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_2_RNI7SOH1_23_LC_9_5_2  (
            .in0(N__3364),
            .in1(N__3097),
            .in2(N__3118),
            .in3(N__3817),
            .lcout(),
            .ltout(\led_blink_inst.o_LED_23_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNIUL825_10_LC_9_5_3 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_RNIUL825_10_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNIUL825_10_LC_9_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_2_RNIUL825_10_LC_9_5_3  (
            .in0(N__2803),
            .in1(N__3178),
            .in2(N__3172),
            .in3(N__3169),
            .lcout(\led_blink_inst.o_LED_23_21 ),
            .ltout(\led_blink_inst.o_LED_23_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_9_LC_9_5_4 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_9_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_9_LC_9_5_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_2_9_LC_9_5_4  (
            .in0(N__3787),
            .in1(N__3723),
            .in2(N__3163),
            .in3(N__3283),
            .lcout(\led_blink_inst.r_Count_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4941),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_4_LC_9_5_5 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_4_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_4_LC_9_5_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_2_4_LC_9_5_5  (
            .in0(N__3722),
            .in1(N__3786),
            .in2(N__3669),
            .in3(N__3070),
            .lcout(\led_blink_inst.r_Count_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4941),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_0_LC_9_5_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_0_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_0_LC_9_5_6 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \led_blink_inst.r_Count_2_0_LC_9_5_6  (
            .in0(N__3137),
            .in1(N__3721),
            .in2(N__3801),
            .in3(N__3646),
            .lcout(\led_blink_inst.r_Count_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4941),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNI3OOH1_21_LC_9_5_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_RNI3OOH1_21_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNI3OOH1_21_LC_9_5_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_2_RNI3OOH1_21_LC_9_5_7  (
            .in0(N__3333),
            .in1(N__3136),
            .in2(N__3847),
            .in3(N__3159),
            .lcout(\led_blink_inst.o_LED_23_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.un2_r_Count_2_1_cry_1_c_LC_9_6_0 .C_ON=1'b1;
    defparam \led_blink_inst.un2_r_Count_2_1_cry_1_c_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.un2_r_Count_2_1_cry_1_c_LC_9_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \led_blink_inst.un2_r_Count_2_1_cry_1_c_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__3153),
            .in2(N__3141),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_2_LC_9_6_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_2_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_2_LC_9_6_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_2_2_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3117),
            .in3(N__3100),
            .lcout(\led_blink_inst.r_Count_2Z0Z_2 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_1 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_2 ),
            .clk(N__4938),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_3_LC_9_6_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_3_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_3_LC_9_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_3_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__3096),
            .in2(_gnd_net_),
            .in3(N__3085),
            .lcout(\led_blink_inst.r_Count_2Z0Z_3 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_2 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_3 ),
            .clk(N__4938),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_4_LC_9_6_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_4_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_4_LC_9_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_4_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__3081),
            .in2(_gnd_net_),
            .in3(N__3064),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_3 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_5_LC_9_6_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_5_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_5_LC_9_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_5_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__3363),
            .in2(_gnd_net_),
            .in3(N__3352),
            .lcout(\led_blink_inst.r_Count_2Z0Z_5 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_4 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_5 ),
            .clk(N__4938),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_6_LC_9_6_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_6_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_6_LC_9_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_6_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(N__3348),
            .in2(_gnd_net_),
            .in3(N__3337),
            .lcout(\led_blink_inst.r_Count_2Z0Z_6 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_5 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_6 ),
            .clk(N__4938),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_7_LC_9_6_6 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_7_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_7_LC_9_6_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_2_7_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3334),
            .in3(N__3319),
            .lcout(\led_blink_inst.r_Count_2Z0Z_7 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_6 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_7 ),
            .clk(N__4938),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_8_LC_9_6_7 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_8_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_8_LC_9_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_8_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__3315),
            .in2(_gnd_net_),
            .in3(N__3304),
            .lcout(\led_blink_inst.r_Count_2Z0Z_8 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_7 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_8 ),
            .clk(N__4938),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_9_LC_9_7_0 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_9_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_9_LC_9_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_9_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__3300),
            .in2(_gnd_net_),
            .in3(N__3274),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_10_LC_9_7_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_10_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_10_LC_9_7_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_10_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3271),
            .in3(N__3247),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_9 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_11_LC_9_7_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_11_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_11_LC_9_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_11_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__3243),
            .in2(_gnd_net_),
            .in3(N__3214),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_10 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_12_LC_9_7_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_12_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_12_LC_9_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_12_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__3210),
            .in2(_gnd_net_),
            .in3(N__3181),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_11 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_13_LC_9_7_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_13_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_13_LC_9_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_13_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__3576),
            .in2(_gnd_net_),
            .in3(N__3565),
            .lcout(\led_blink_inst.r_Count_2Z0Z_13 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_12 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_13 ),
            .clk(N__4935),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_14_LC_9_7_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_14_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_14_LC_9_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_14_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__3561),
            .in2(_gnd_net_),
            .in3(N__3544),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_13 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_15_LC_9_7_6 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_15_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_15_LC_9_7_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_2_15_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3540),
            .in3(N__3523),
            .lcout(\led_blink_inst.r_Count_2Z0Z_15 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_14 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_15 ),
            .clk(N__4935),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_16_LC_9_7_7 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_16_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_16_LC_9_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_16_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__3520),
            .in2(_gnd_net_),
            .in3(N__3496),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_15 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_17_LC_9_8_0 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_17_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_17_LC_9_8_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_17_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3493),
            .in3(N__3460),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_18_LC_9_8_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_18_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_18_LC_9_8_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_18_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3457),
            .in3(N__3430),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_17 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_19_LC_9_8_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_19_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_19_LC_9_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_19_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__3427),
            .in2(_gnd_net_),
            .in3(N__3400),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_18 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_20_LC_9_8_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_20_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_20_LC_9_8_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_20_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3397),
            .in3(N__3367),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_19 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_21_LC_9_8_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_21_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_21_LC_9_8_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_2_21_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3843),
            .in3(N__3826),
            .lcout(\led_blink_inst.r_Count_2Z0Z_21 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_20 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_21 ),
            .clk(N__4931),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_RNO_0_22_LC_9_8_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_2_RNO_0_22_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_2_RNO_0_22_LC_9_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_2_RNO_0_22_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__3594),
            .in2(_gnd_net_),
            .in3(N__3823),
            .lcout(\led_blink_inst.r_Count_2_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_2_1_cry_21 ),
            .carryout(\led_blink_inst.un2_r_Count_2_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_23_LC_9_8_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_23_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_23_LC_9_8_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \led_blink_inst.r_Count_2_23_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__3816),
            .in2(_gnd_net_),
            .in3(N__3820),
            .lcout(\led_blink_inst.r_Count_2Z0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4931),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_2_22_LC_9_8_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_2_22_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_2_22_LC_9_8_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_2_22_LC_9_8_7  (
            .in0(N__3802),
            .in1(N__3739),
            .in2(N__3682),
            .in3(N__3673),
            .lcout(\led_blink_inst.r_Count_2Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4931),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNI527P1_11_LC_11_3_1 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_RNI527P1_11_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNI527P1_11_LC_11_3_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_3_RNI527P1_11_LC_11_3_1  (
            .in0(N__4297),
            .in1(N__4113),
            .in2(N__4435),
            .in3(N__4266),
            .lcout(\led_blink_inst.o_LED_33_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_8_LC_11_3_2 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_8_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_8_LC_11_3_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_3_8_LC_11_3_2  (
            .in0(N__4038),
            .in1(N__3994),
            .in2(N__4171),
            .in3(N__3954),
            .lcout(\led_blink_inst.r_Count_3Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4949),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_7_LC_11_3_4 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_7_LC_11_3_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_7_LC_11_3_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_3_7_LC_11_3_4  (
            .in0(N__4037),
            .in1(N__3993),
            .in2(N__3958),
            .in3(N__4195),
            .lcout(\led_blink_inst.r_Count_3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4949),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNIHE7P1_10_LC_11_3_5 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_RNIHE7P1_10_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNIHE7P1_10_LC_11_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_3_RNIHE7P1_10_LC_11_3_5  (
            .in0(N__4210),
            .in1(N__4249),
            .in2(N__4462),
            .in3(N__4185),
            .lcout(\led_blink_inst.o_LED_33_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_5_LC_11_3_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_5_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_5_LC_11_3_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_3_5_LC_11_3_6  (
            .in0(N__4036),
            .in1(N__3992),
            .in2(N__3957),
            .in3(N__4237),
            .lcout(\led_blink_inst.r_Count_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4949),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_1_LC_11_3_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_1_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_1_LC_11_3_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_1_LC_11_3_7  (
            .in0(N__4098),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4114),
            .lcout(\led_blink_inst.r_Count_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4949),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNIU40L1_23_LC_11_4_0 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_RNIU40L1_23_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNIU40L1_23_LC_11_4_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_3_RNIU40L1_23_LC_11_4_0  (
            .in0(N__4338),
            .in1(N__4228),
            .in2(N__4507),
            .in3(N__4096),
            .lcout(\led_blink_inst.o_LED_33_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNIK2NG1_14_LC_11_4_1 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_RNIK2NG1_14_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNIK2NG1_14_LC_11_4_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_3_RNIK2NG1_14_LC_11_4_1  (
            .in0(N__4375),
            .in1(N__4282),
            .in2(N__4591),
            .in3(N__4356),
            .lcout(),
            .ltout(\led_blink_inst.o_LED_33_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNIEFLF6_10_LC_11_4_2 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_RNIEFLF6_10_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNIEFLF6_10_LC_11_4_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_3_RNIEFLF6_10_LC_11_4_2  (
            .in0(N__3892),
            .in1(N__3883),
            .in2(N__3877),
            .in3(N__4048),
            .lcout(\led_blink_inst.o_LED_33_21 ),
            .ltout(\led_blink_inst.o_LED_33_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.o_LED_3_LC_11_4_3 .C_ON=1'b0;
    defparam \led_blink_inst.o_LED_3_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.o_LED_3_LC_11_4_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \led_blink_inst.o_LED_3_LC_11_4_3  (
            .in0(N__3867),
            .in1(N__4023),
            .in2(N__3874),
            .in3(N__3986),
            .lcout(o_LED_3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4947),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_10_LC_11_4_4 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_10_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_10_LC_11_4_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_3_10_LC_11_4_4  (
            .in0(N__3988),
            .in1(N__4027),
            .in2(N__3955),
            .in3(N__4444),
            .lcout(\led_blink_inst.r_Count_3Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4947),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNIEUOG1_12_LC_11_4_5 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_RNIEUOG1_12_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNIEUOG1_12_LC_11_4_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_3_RNIEUOG1_12_LC_11_4_5  (
            .in0(N__4569),
            .in1(N__4413),
            .in2(N__4528),
            .in3(N__4155),
            .lcout(\led_blink_inst.o_LED_33_16 ),
            .ltout(\led_blink_inst.o_LED_33_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_13_LC_11_4_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_13_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_13_LC_11_4_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_3_13_LC_11_4_6  (
            .in0(N__3941),
            .in1(N__4028),
            .in2(N__3850),
            .in3(N__4384),
            .lcout(\led_blink_inst.r_Count_3Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4947),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_0_LC_11_4_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_0_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_0_LC_11_4_7 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \led_blink_inst.r_Count_3_0_LC_11_4_7  (
            .in0(N__4097),
            .in1(N__3987),
            .in2(N__4039),
            .in3(N__3942),
            .lcout(\led_blink_inst.r_Count_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4947),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_21_LC_11_5_0 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_21_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_21_LC_11_5_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_3_21_LC_11_5_0  (
            .in0(N__3991),
            .in1(N__4042),
            .in2(N__3956),
            .in3(N__4537),
            .lcout(\led_blink_inst.r_Count_3Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4945),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_17_LC_11_5_1 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_17_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_17_LC_11_5_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_3_17_LC_11_5_1  (
            .in0(N__4040),
            .in1(N__3989),
            .in2(N__4309),
            .in3(N__3946),
            .lcout(\led_blink_inst.r_Count_3Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4945),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNI4SFC1_13_LC_11_5_3 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_RNI4SFC1_13_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNI4SFC1_13_LC_11_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_3_RNI4SFC1_13_LC_11_5_3  (
            .in0(N__4320),
            .in1(N__4396),
            .in2(N__4552),
            .in3(N__4617),
            .lcout(\led_blink_inst.o_LED_33_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_18_LC_11_5_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_18_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_18_LC_11_5_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_3_18_LC_11_5_7  (
            .in0(N__4041),
            .in1(N__3990),
            .in2(N__4603),
            .in3(N__3947),
            .lcout(\led_blink_inst.r_Count_3Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4945),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.un2_r_Count_4_1_cry_1_c_LC_11_6_0 .C_ON=1'b1;
    defparam \led_blink_inst.un2_r_Count_4_1_cry_1_c_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.un2_r_Count_4_1_cry_1_c_LC_11_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \led_blink_inst.un2_r_Count_4_1_cry_1_c_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__5170),
            .in2(N__5136),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_2_LC_11_6_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_2_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_2_LC_11_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_2_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__5244),
            .in2(_gnd_net_),
            .in3(N__3907),
            .lcout(\led_blink_inst.r_Count_4Z0Z_2 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_1 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_2 ),
            .clk(N__4942),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_3_LC_11_6_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_3_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_3_LC_11_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_3_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__4629),
            .in2(_gnd_net_),
            .in3(N__3904),
            .lcout(\led_blink_inst.r_Count_4Z0Z_3 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_2 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_3 ),
            .clk(N__4942),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNO_0_4_LC_11_6_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_RNO_0_4_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNO_0_4_LC_11_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_RNO_0_4_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__4761),
            .in2(_gnd_net_),
            .in3(N__3901),
            .lcout(\led_blink_inst.r_Count_4_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_3 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_5_LC_11_6_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_5_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_5_LC_11_6_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_4_5_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4705),
            .in3(N__3898),
            .lcout(\led_blink_inst.r_Count_4Z0Z_5 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_4 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_5 ),
            .clk(N__4942),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNO_0_6_LC_11_6_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_RNO_0_6_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNO_0_6_LC_11_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_RNO_0_6_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__4800),
            .in2(_gnd_net_),
            .in3(N__3895),
            .lcout(\led_blink_inst.r_Count_4_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_5 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNO_0_7_LC_11_6_6 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_RNO_0_7_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNO_0_7_LC_11_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_RNO_0_7_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(N__4773),
            .in2(_gnd_net_),
            .in3(N__4075),
            .lcout(\led_blink_inst.r_Count_4_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_6 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_8_LC_11_6_7 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_8_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_8_LC_11_6_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_4_8_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4750),
            .in3(N__4072),
            .lcout(\led_blink_inst.r_Count_4Z0Z_8 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_7 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_8 ),
            .clk(N__4942),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNO_0_9_LC_11_7_0 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_RNO_0_9_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNO_0_9_LC_11_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_RNO_0_9_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__4788),
            .in2(_gnd_net_),
            .in3(N__4069),
            .lcout(\led_blink_inst.r_Count_4_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_10_LC_11_7_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_10_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_10_LC_11_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_10_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__4734),
            .in2(_gnd_net_),
            .in3(N__4066),
            .lcout(\led_blink_inst.r_Count_4Z0Z_10 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_9 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_10 ),
            .clk(N__4940),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_11_LC_11_7_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_11_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_11_LC_11_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_11_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__5256),
            .in2(_gnd_net_),
            .in3(N__4063),
            .lcout(\led_blink_inst.r_Count_4Z0Z_11 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_10 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_11 ),
            .clk(N__4940),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNO_0_12_LC_11_7_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_RNO_0_12_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNO_0_12_LC_11_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_RNO_0_12_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__4870),
            .in2(_gnd_net_),
            .in3(N__4060),
            .lcout(\led_blink_inst.r_Count_4_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_11 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_13_LC_11_7_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_13_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_13_LC_11_7_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_4_13_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4722),
            .in3(N__4057),
            .lcout(\led_blink_inst.r_Count_4Z0Z_13 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_12 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_13 ),
            .clk(N__4940),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_14_LC_11_7_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_14_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_14_LC_11_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_14_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__4668),
            .in2(_gnd_net_),
            .in3(N__4054),
            .lcout(\led_blink_inst.r_Count_4Z0Z_14 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_13 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_14 ),
            .clk(N__4940),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_15_LC_11_7_6 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_15_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_15_LC_11_7_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_4_15_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5215),
            .in3(N__4051),
            .lcout(\led_blink_inst.r_Count_4Z0Z_15 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_14 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_15 ),
            .clk(N__4940),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNO_0_16_LC_11_7_7 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_RNO_0_16_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNO_0_16_LC_11_7_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_4_RNO_0_16_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4855),
            .in3(N__4138),
            .lcout(\led_blink_inst.r_Count_4_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_15 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNO_0_17_LC_11_8_0 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_RNO_0_17_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNO_0_17_LC_11_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_RNO_0_17_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__4839),
            .in2(_gnd_net_),
            .in3(N__4135),
            .lcout(\led_blink_inst.r_Count_4_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_18_LC_11_8_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_18_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_18_LC_11_8_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_4_18_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5232),
            .in3(N__4132),
            .lcout(\led_blink_inst.r_Count_4Z0Z_18 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_17 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_18 ),
            .clk(N__4936),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_19_LC_11_8_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_19_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_19_LC_11_8_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_4_19_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5191),
            .in3(N__4129),
            .lcout(\led_blink_inst.r_Count_4Z0Z_19 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_18 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_19 ),
            .clk(N__4936),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNO_0_20_LC_11_8_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_RNO_0_20_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNO_0_20_LC_11_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_RNO_0_20_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__4825),
            .in2(_gnd_net_),
            .in3(N__4126),
            .lcout(\led_blink_inst.r_Count_4_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_19 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_21_LC_11_8_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_21_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_21_LC_11_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_21_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__4644),
            .in2(_gnd_net_),
            .in3(N__4123),
            .lcout(\led_blink_inst.r_Count_4Z0Z_21 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_20 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_21 ),
            .clk(N__4936),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_22_LC_11_8_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_4_22_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_22_LC_11_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_4_22_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__5151),
            .in2(_gnd_net_),
            .in3(N__4120),
            .lcout(\led_blink_inst.r_Count_4Z0Z_22 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_4_1_cry_21 ),
            .carryout(\led_blink_inst.un2_r_Count_4_1_cry_22 ),
            .clk(N__4936),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_23_LC_11_8_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_23_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_23_LC_11_8_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \led_blink_inst.r_Count_4_23_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__4657),
            .in2(_gnd_net_),
            .in3(N__4117),
            .lcout(\led_blink_inst.r_Count_4Z0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4936),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.un2_r_Count_3_1_cry_1_c_LC_12_3_0 .C_ON=1'b1;
    defparam \led_blink_inst.un2_r_Count_3_1_cry_1_c_LC_12_3_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.un2_r_Count_3_1_cry_1_c_LC_12_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \led_blink_inst.un2_r_Count_3_1_cry_1_c_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(N__4112),
            .in2(N__4099),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_3_0_),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_2_LC_12_3_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_2_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_2_LC_12_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_3_2_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(N__4296),
            .in2(_gnd_net_),
            .in3(N__4285),
            .lcout(\led_blink_inst.r_Count_3Z0Z_2 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_1 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_2 ),
            .clk(N__4951),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_3_LC_12_3_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_3_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_3_LC_12_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_3_3_LC_12_3_2  (
            .in0(_gnd_net_),
            .in1(N__4281),
            .in2(_gnd_net_),
            .in3(N__4270),
            .lcout(\led_blink_inst.r_Count_3Z0Z_3 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_2 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_3 ),
            .clk(N__4951),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_4_LC_12_3_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_4_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_4_LC_12_3_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_4_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4267),
            .in3(N__4252),
            .lcout(\led_blink_inst.r_Count_3Z0Z_4 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_3 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_4 ),
            .clk(N__4951),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNO_0_5_LC_12_3_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_RNO_0_5_LC_12_3_4 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNO_0_5_LC_12_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_3_RNO_0_5_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(N__4248),
            .in2(_gnd_net_),
            .in3(N__4231),
            .lcout(\led_blink_inst.r_Count_3_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_4 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_6_LC_12_3_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_6_LC_12_3_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_6_LC_12_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_3_6_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(N__4224),
            .in2(_gnd_net_),
            .in3(N__4213),
            .lcout(\led_blink_inst.r_Count_3Z0Z_6 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_5 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_6 ),
            .clk(N__4951),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNO_0_7_LC_12_3_6 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_RNO_0_7_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNO_0_7_LC_12_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_3_RNO_0_7_LC_12_3_6  (
            .in0(_gnd_net_),
            .in1(N__4206),
            .in2(_gnd_net_),
            .in3(N__4189),
            .lcout(\led_blink_inst.r_Count_3_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_6 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNO_0_8_LC_12_3_7 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_RNO_0_8_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNO_0_8_LC_12_3_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_RNO_0_8_LC_12_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4186),
            .in3(N__4159),
            .lcout(\led_blink_inst.r_Count_3_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_7 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_9_LC_12_4_0 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_9_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_9_LC_12_4_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_9_LC_12_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4156),
            .in3(N__4141),
            .lcout(\led_blink_inst.r_Count_3Z0Z_9 ),
            .ltout(),
            .carryin(bfn_12_4_0_),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_9 ),
            .clk(N__4950),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNO_0_10_LC_12_4_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_RNO_0_10_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNO_0_10_LC_12_4_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_RNO_0_10_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4461),
            .in3(N__4438),
            .lcout(\led_blink_inst.r_Count_3_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_9 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_11_LC_12_4_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_11_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_11_LC_12_4_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_11_LC_12_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4434),
            .in3(N__4417),
            .lcout(\led_blink_inst.r_Count_3Z0Z_11 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_10 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_11 ),
            .clk(N__4950),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_12_LC_12_4_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_12_LC_12_4_3 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_12_LC_12_4_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_12_LC_12_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4414),
            .in3(N__4399),
            .lcout(\led_blink_inst.r_Count_3Z0Z_12 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_11 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_12 ),
            .clk(N__4950),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNO_0_13_LC_12_4_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_RNO_0_13_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNO_0_13_LC_12_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_3_RNO_0_13_LC_12_4_4  (
            .in0(_gnd_net_),
            .in1(N__4395),
            .in2(_gnd_net_),
            .in3(N__4378),
            .lcout(\led_blink_inst.r_Count_3_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_12 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_14_LC_12_4_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_14_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_14_LC_12_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_3_14_LC_12_4_5  (
            .in0(_gnd_net_),
            .in1(N__4371),
            .in2(_gnd_net_),
            .in3(N__4360),
            .lcout(\led_blink_inst.r_Count_3Z0Z_14 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_13 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_14 ),
            .clk(N__4950),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_15_LC_12_4_6 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_15_LC_12_4_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_15_LC_12_4_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_15_LC_12_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4357),
            .in3(N__4342),
            .lcout(\led_blink_inst.r_Count_3Z0Z_15 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_14 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_15 ),
            .clk(N__4950),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_16_LC_12_4_7 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_16_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_16_LC_12_4_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_16_LC_12_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4339),
            .in3(N__4324),
            .lcout(\led_blink_inst.r_Count_3Z0Z_16 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_15 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_16 ),
            .clk(N__4950),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNO_0_17_LC_12_5_0 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_RNO_0_17_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNO_0_17_LC_12_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_3_RNO_0_17_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__4321),
            .in2(_gnd_net_),
            .in3(N__4300),
            .lcout(\led_blink_inst.r_Count_3_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNO_0_18_LC_12_5_1 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_RNO_0_18_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNO_0_18_LC_12_5_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_RNO_0_18_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4618),
            .in3(N__4594),
            .lcout(\led_blink_inst.r_Count_3_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_17 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_19_LC_12_5_2 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_19_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_19_LC_12_5_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_19_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4590),
            .in3(N__4573),
            .lcout(\led_blink_inst.r_Count_3Z0Z_19 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_18 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_19 ),
            .clk(N__4948),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_20_LC_12_5_3 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_20_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_20_LC_12_5_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_3_20_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4570),
            .in3(N__4555),
            .lcout(\led_blink_inst.r_Count_3Z0Z_20 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_19 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_20 ),
            .clk(N__4948),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_RNO_0_21_LC_12_5_4 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_RNO_0_21_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_3_RNO_0_21_LC_12_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_3_RNO_0_21_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(N__4551),
            .in2(_gnd_net_),
            .in3(N__4531),
            .lcout(\led_blink_inst.r_Count_3_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_20 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_22_LC_12_5_5 .C_ON=1'b1;
    defparam \led_blink_inst.r_Count_3_22_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_22_LC_12_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \led_blink_inst.r_Count_3_22_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(N__4527),
            .in2(_gnd_net_),
            .in3(N__4513),
            .lcout(\led_blink_inst.r_Count_3Z0Z_22 ),
            .ltout(),
            .carryin(\led_blink_inst.un2_r_Count_3_1_cry_21 ),
            .carryout(\led_blink_inst.un2_r_Count_3_1_cry_22 ),
            .clk(N__4948),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_3_23_LC_12_5_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_3_23_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_3_23_LC_12_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \led_blink_inst.r_Count_3_23_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(N__4503),
            .in2(_gnd_net_),
            .in3(N__4510),
            .lcout(\led_blink_inst.r_Count_3Z0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4948),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_4_LC_12_6_0 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_4_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_4_LC_12_6_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_4_4_LC_12_6_0  (
            .in0(N__4992),
            .in1(N__5037),
            .in2(N__4489),
            .in3(N__5087),
            .lcout(\led_blink_inst.r_Count_4Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4946),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_7_LC_12_6_1 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_7_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_7_LC_12_6_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_4_7_LC_12_6_1  (
            .in0(N__5039),
            .in1(N__4989),
            .in2(N__5091),
            .in3(N__4477),
            .lcout(\led_blink_inst.r_Count_4Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4946),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_6_LC_12_6_2 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_6_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_6_LC_12_6_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_4_6_LC_12_6_2  (
            .in0(N__4993),
            .in1(N__5038),
            .in2(N__4471),
            .in3(N__5088),
            .lcout(\led_blink_inst.r_Count_4Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4946),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_9_LC_12_6_3 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_9_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_9_LC_12_6_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_4_9_LC_12_6_3  (
            .in0(N__5040),
            .in1(N__4990),
            .in2(N__5092),
            .in3(N__4807),
            .lcout(\led_blink_inst.r_Count_4Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4946),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNIA7S1_4_LC_12_6_4 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_RNIA7S1_4_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNIA7S1_4_LC_12_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_4_RNIA7S1_4_LC_12_6_4  (
            .in0(N__4801),
            .in1(N__4789),
            .in2(N__4777),
            .in3(N__4762),
            .lcout(\led_blink_inst.o_LED_43_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNI2IHV_5_LC_12_6_5 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_RNI2IHV_5_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNI2IHV_5_LC_12_6_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_4_RNI2IHV_5_LC_12_6_5  (
            .in0(N__4749),
            .in1(N__4735),
            .in2(N__4723),
            .in3(N__4704),
            .lcout(\led_blink_inst.o_LED_43_16 ),
            .ltout(\led_blink_inst.o_LED_43_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_0_LC_12_6_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_0_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_0_LC_12_6_6 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \led_blink_inst.r_Count_4_0_LC_12_6_6  (
            .in0(N__4991),
            .in1(N__5086),
            .in2(N__4690),
            .in3(N__5174),
            .lcout(\led_blink_inst.r_Count_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4946),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_1_LC_12_6_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_1_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_1_LC_12_6_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \led_blink_inst.r_Count_4_1_LC_12_6_7  (
            .in0(N__5175),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5135),
            .lcout(\led_blink_inst.r_Count_4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4946),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_16_LC_12_7_0 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_16_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_16_LC_12_7_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_4_16_LC_12_7_0  (
            .in0(N__5036),
            .in1(N__5090),
            .in2(N__4994),
            .in3(N__4687),
            .lcout(\led_blink_inst.r_Count_4Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4943),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_12_LC_12_7_1 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_12_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_12_LC_12_7_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_4_12_LC_12_7_1  (
            .in0(N__5089),
            .in1(N__5035),
            .in2(N__4681),
            .in3(N__4983),
            .lcout(\led_blink_inst.r_Count_4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4943),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNIGBEE1_23_LC_12_7_2 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_RNIGBEE1_23_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNIGBEE1_23_LC_12_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_4_RNIGBEE1_23_LC_12_7_2  (
            .in0(N__4672),
            .in1(N__4656),
            .in2(N__4645),
            .in3(N__4630),
            .lcout(),
            .ltout(\led_blink_inst.o_LED_43_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNIH7VR4_2_LC_12_7_3 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_RNIH7VR4_2_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNIH7VR4_2_LC_12_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_4_RNIH7VR4_2_LC_12_7_3  (
            .in0(N__5200),
            .in1(N__4813),
            .in2(N__5266),
            .in3(N__5263),
            .lcout(\led_blink_inst.o_LED_43_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNIJCCE1_2_LC_12_7_4 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_RNIJCCE1_2_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNIJCCE1_2_LC_12_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_4_RNIJCCE1_2_LC_12_7_4  (
            .in0(N__5257),
            .in1(N__5245),
            .in2(N__5233),
            .in3(N__5214),
            .lcout(\led_blink_inst.o_LED_43_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNIVFIV_1_LC_12_7_6 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_RNIVFIV_1_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNIVFIV_1_LC_12_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \led_blink_inst.r_Count_4_RNIVFIV_1_LC_12_7_6  (
            .in0(N__5190),
            .in1(N__5176),
            .in2(N__5152),
            .in3(N__5137),
            .lcout(\led_blink_inst.o_LED_43_17 ),
            .ltout(\led_blink_inst.o_LED_43_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.o_LED_4_LC_12_7_7 .C_ON=1'b0;
    defparam \led_blink_inst.o_LED_4_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.o_LED_4_LC_12_7_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \led_blink_inst.o_LED_4_LC_12_7_7  (
            .in0(N__5109),
            .in1(N__5034),
            .in2(N__5113),
            .in3(N__4982),
            .lcout(o_LED_4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4943),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_20_LC_12_8_0 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_20_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_20_LC_12_8_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \led_blink_inst.r_Count_4_20_LC_12_8_0  (
            .in0(N__5047),
            .in1(N__5079),
            .in2(N__4999),
            .in3(N__5098),
            .lcout(\led_blink_inst.r_Count_4Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4939),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_17_LC_12_8_3 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_17_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \led_blink_inst.r_Count_4_17_LC_12_8_3 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \led_blink_inst.r_Count_4_17_LC_12_8_3  (
            .in0(N__5078),
            .in1(N__5046),
            .in2(N__5008),
            .in3(N__4998),
            .lcout(\led_blink_inst.r_Count_4Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4939),
            .ce(),
            .sr(_gnd_net_));
    defparam \led_blink_inst.r_Count_4_RNI488T1_12_LC_12_8_7 .C_ON=1'b0;
    defparam \led_blink_inst.r_Count_4_RNI488T1_12_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \led_blink_inst.r_Count_4_RNI488T1_12_LC_12_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \led_blink_inst.r_Count_4_RNI488T1_12_LC_12_8_7  (
            .in0(N__4869),
            .in1(N__4854),
            .in2(N__4840),
            .in3(N__4824),
            .lcout(\led_blink_inst.o_LED_43_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // led_blink_top
