module hello_world_tb();
  
  // due to initial block, the messgae is displayed only once
  initial $display("Hello, World!");
  
endmodule
