-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jul 24 2022 20:50:09

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "led_blink_top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of led_blink_top
entity led_blink_top is
port (
    o_LED_3 : out std_logic;
    o_LED_1 : out std_logic;
    i_Clk : in std_logic;
    o_LED_4 : out std_logic;
    o_LED_2 : out std_logic);
end led_blink_top;

-- Architecture of led_blink_top
-- View name is \INTERFACE\
architecture \INTERFACE\ of led_blink_top is

signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2527\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2359\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2302\ : std_logic;
signal \N__2299\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2293\ : std_logic;
signal \N__2290\ : std_logic;
signal \N__2287\ : std_logic;
signal \N__2284\ : std_logic;
signal \N__2281\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2259\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \o_LED_1_c\ : std_logic;
signal \led_blink_inst.o_LED_13_15\ : std_logic;
signal \led_blink_inst.o_LED_13_13\ : std_logic;
signal \led_blink_inst.o_LED_13_14_cascade_\ : std_logic;
signal \led_blink_inst.o_LED_13_12\ : std_logic;
signal \led_blink_inst.o_LED_13_21_cascade_\ : std_logic;
signal \led_blink_inst.o_LED_13_16_cascade_\ : std_logic;
signal \led_blink_inst.o_LED_23_16_cascade_\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_1\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_0\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_2\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_1\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_3\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_2\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_4\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_3\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_5\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_5\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_4\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_6\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_5\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_7\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_6\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_8\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_7\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_8\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_9\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_10\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_10\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_9\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_11\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_11\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_10\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_12\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_12\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_11\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_13\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_13\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_12\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_14\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_13\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_15\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_15\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_14\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_16\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_15\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_16\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_17\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_17\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_18\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_18\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_17\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_19\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_19\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_18\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_20\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_20\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_19\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_21\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_21\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_20\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_22\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_21\ : std_logic;
signal \led_blink_inst.un3_r_Count_1_1_cry_22\ : std_logic;
signal \led_blink_inst.o_LED_13_17\ : std_logic;
signal \led_blink_inst.o_LED_13_16\ : std_logic;
signal \led_blink_inst.r_Count_1_RNO_0Z0Z_23_cascade_\ : std_logic;
signal \led_blink_inst.o_LED_13_21\ : std_logic;
signal \led_blink_inst.r_Count_1Z0Z_23\ : std_logic;
signal \o_LED_2_c\ : std_logic;
signal \led_blink_inst.o_LED_23_14\ : std_logic;
signal \led_blink_inst.o_LED_23_13\ : std_logic;
signal \led_blink_inst.o_LED_23_12_cascade_\ : std_logic;
signal \led_blink_inst.o_LED_23_15\ : std_logic;
signal \led_blink_inst.o_LED_23_21_cascade_\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_1\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_0\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_2\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_1\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_3\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_2\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_4\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_4\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_3\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_5\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_4\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_6\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_5\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_7\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_6\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_8\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_7\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_8\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_9\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_9\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_10\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_10\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_9\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_11\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_11\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_10\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_12\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_12\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_11\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_13\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_12\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_14\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_14\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_13\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_15\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_14\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_16\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_16\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_15\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_16\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_17\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_17\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_18\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_18\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_17\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_19\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_19\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_18\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_20\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_20\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_19\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_21\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_20\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_21\ : std_logic;
signal \led_blink_inst.un2_r_Count_2_1_cry_22\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_23\ : std_logic;
signal \led_blink_inst.o_LED_23_17\ : std_logic;
signal \led_blink_inst.o_LED_23_16\ : std_logic;
signal \led_blink_inst.r_Count_2_RNO_0Z0Z_22\ : std_logic;
signal \led_blink_inst.o_LED_23_21\ : std_logic;
signal \led_blink_inst.r_Count_2Z0Z_22\ : std_logic;
signal \led_blink_inst.o_LED_33_14\ : std_logic;
signal \led_blink_inst.o_LED_33_13\ : std_logic;
signal \led_blink_inst.o_LED_33_12_cascade_\ : std_logic;
signal \led_blink_inst.o_LED_33_21_cascade_\ : std_logic;
signal \o_LED_3_c\ : std_logic;
signal \led_blink_inst.o_LED_33_16_cascade_\ : std_logic;
signal \led_blink_inst.o_LED_33_15\ : std_logic;
signal \led_blink_inst.o_LED_33_17\ : std_logic;
signal \led_blink_inst.o_LED_33_16\ : std_logic;
signal \led_blink_inst.o_LED_33_21\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_1\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_2\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_3\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_4\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_5\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_6\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_7\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_8\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_9\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_10\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_11\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_12\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_13\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_14\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_15\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_16\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_17\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_18\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_19\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_20\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_21\ : std_logic;
signal \led_blink_inst.un2_r_Count_4_1_cry_22\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_1\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_0\ : std_logic;
signal \bfn_12_3_0_\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_2\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_1\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_3\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_2\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_4\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_3\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_5\ : std_logic;
signal \led_blink_inst.r_Count_3_RNO_0Z0Z_5\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_4\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_6\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_5\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_7\ : std_logic;
signal \led_blink_inst.r_Count_3_RNO_0Z0Z_7\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_6\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_8\ : std_logic;
signal \led_blink_inst.r_Count_3_RNO_0Z0Z_8\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_7\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_8\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_9\ : std_logic;
signal \bfn_12_4_0_\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_10\ : std_logic;
signal \led_blink_inst.r_Count_3_RNO_0Z0Z_10\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_9\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_11\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_10\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_12\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_11\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_13\ : std_logic;
signal \led_blink_inst.r_Count_3_RNO_0Z0Z_13\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_12\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_14\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_13\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_15\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_14\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_16\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_15\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_16\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_17\ : std_logic;
signal \led_blink_inst.r_Count_3_RNO_0Z0Z_17\ : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_18\ : std_logic;
signal \led_blink_inst.r_Count_3_RNO_0Z0Z_18\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_17\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_19\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_18\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_20\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_19\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_21\ : std_logic;
signal \led_blink_inst.r_Count_3_RNO_0Z0Z_21\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_20\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_22\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_21\ : std_logic;
signal \led_blink_inst.un2_r_Count_3_1_cry_22\ : std_logic;
signal \led_blink_inst.r_Count_3Z0Z_23\ : std_logic;
signal \led_blink_inst.r_Count_4_RNO_0Z0Z_4\ : std_logic;
signal \led_blink_inst.r_Count_4_RNO_0Z0Z_7\ : std_logic;
signal \led_blink_inst.r_Count_4_RNO_0Z0Z_6\ : std_logic;
signal \led_blink_inst.r_Count_4_RNO_0Z0Z_9\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_6\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_9\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_7\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_4\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_8\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_10\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_13\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_5\ : std_logic;
signal \led_blink_inst.o_LED_43_16_cascade_\ : std_logic;
signal \led_blink_inst.r_Count_4_RNO_0Z0Z_16\ : std_logic;
signal \led_blink_inst.r_Count_4_RNO_0Z0Z_12\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_14\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_23\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_21\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_3\ : std_logic;
signal \led_blink_inst.o_LED_43_12_cascade_\ : std_logic;
signal \led_blink_inst.o_LED_43_14\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_11\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_2\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_18\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_15\ : std_logic;
signal \led_blink_inst.o_LED_43_13\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_19\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_0\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_22\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_1\ : std_logic;
signal \led_blink_inst.o_LED_43_17_cascade_\ : std_logic;
signal \o_LED_4_c\ : std_logic;
signal \led_blink_inst.r_Count_4_RNO_0Z0Z_20\ : std_logic;
signal \led_blink_inst.o_LED_43_17\ : std_logic;
signal \led_blink_inst.o_LED_43_16\ : std_logic;
signal \led_blink_inst.r_Count_4_RNO_0Z0Z_17\ : std_logic;
signal \led_blink_inst.o_LED_43_21\ : std_logic;
signal \i_Clk_c_g\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_12\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_16\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_17\ : std_logic;
signal \led_blink_inst.r_Count_4Z0Z_20\ : std_logic;
signal \led_blink_inst.o_LED_43_15\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \i_Clk_wire\ : std_logic;
signal \o_LED_1_wire\ : std_logic;
signal \o_LED_2_wire\ : std_logic;
signal \o_LED_3_wire\ : std_logic;
signal \o_LED_4_wire\ : std_logic;

begin
    \i_Clk_wire\ <= i_Clk;
    o_LED_1 <= \o_LED_1_wire\;
    o_LED_2 <= \o_LED_2_wire\;
    o_LED_3 <= \o_LED_3_wire\;
    o_LED_4 <= \o_LED_4_wire\;

    \i_Clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5321\,
            GLOBALBUFFEROUTPUT => \i_Clk_c_g\
        );

    \i_Clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5323\,
            DIN => \N__5322\,
            DOUT => \N__5321\,
            PACKAGEPIN => \i_Clk_wire\
        );

    \i_Clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5323\,
            PADOUT => \N__5322\,
            PADIN => \N__5321\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5312\,
            DIN => \N__5311\,
            DOUT => \N__5310\,
            PACKAGEPIN => \o_LED_1_wire\
        );

    \o_LED_1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5312\,
            PADOUT => \N__5311\,
            PADIN => \N__5310\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2275\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5303\,
            DIN => \N__5302\,
            DOUT => \N__5301\,
            PACKAGEPIN => \o_LED_2_wire\
        );

    \o_LED_2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5303\,
            PADOUT => \N__5302\,
            PADIN => \N__5301\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2824\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5294\,
            DIN => \N__5293\,
            DOUT => \N__5292\,
            PACKAGEPIN => \o_LED_3_wire\
        );

    \o_LED_3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5294\,
            PADOUT => \N__5293\,
            PADIN => \N__5292\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3871\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5285\,
            DIN => \N__5284\,
            DOUT => \N__5283\,
            PACKAGEPIN => \o_LED_4_wire\
        );

    \o_LED_4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5285\,
            PADOUT => \N__5284\,
            PADIN => \N__5283\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5110\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__5266\,
            I => \led_blink_inst.o_LED_43_12_cascade_\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5260\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5260\,
            I => \led_blink_inst.o_LED_43_14\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5253\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5250\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5253\,
            I => \led_blink_inst.r_Count_4Z0Z_11\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5250\,
            I => \led_blink_inst.r_Count_4Z0Z_11\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5245\,
            I => \N__5241\
        );

    \I__1187\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5238\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5241\,
            I => \led_blink_inst.r_Count_4Z0Z_2\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5238\,
            I => \led_blink_inst.r_Count_4Z0Z_2\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__5233\,
            I => \N__5229\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__5232\,
            I => \N__5226\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5223\
        );

    \I__1181\ : InMux
    port map (
            O => \N__5226\,
            I => \N__5220\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5223\,
            I => \led_blink_inst.r_Count_4Z0Z_18\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5220\,
            I => \led_blink_inst.r_Count_4Z0Z_18\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__5215\,
            I => \N__5211\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5208\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5205\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__5208\,
            I => \led_blink_inst.r_Count_4Z0Z_15\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__5205\,
            I => \led_blink_inst.r_Count_4Z0Z_15\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5197\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__5197\,
            I => \N__5194\
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__5194\,
            I => \led_blink_inst.o_LED_43_13\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__5191\,
            I => \N__5187\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5190\,
            I => \N__5184\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5181\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5184\,
            I => \led_blink_inst.r_Count_4Z0Z_19\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5181\,
            I => \led_blink_inst.r_Count_4Z0Z_19\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5171\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5175\,
            I => \N__5165\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5174\,
            I => \N__5165\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__5171\,
            I => \N__5162\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5159\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5165\,
            I => \led_blink_inst.r_Count_4Z0Z_0\
        );

    \I__1159\ : Odrv4
    port map (
            O => \N__5162\,
            I => \led_blink_inst.r_Count_4Z0Z_0\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5159\,
            I => \led_blink_inst.r_Count_4Z0Z_0\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__5152\,
            I => \N__5148\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5145\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5142\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5145\,
            I => \led_blink_inst.r_Count_4Z0Z_22\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5142\,
            I => \led_blink_inst.r_Count_4Z0Z_22\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5132\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__5136\,
            I => \N__5129\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5135\,
            I => \N__5126\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5132\,
            I => \N__5123\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5120\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5126\,
            I => \led_blink_inst.r_Count_4Z0Z_1\
        );

    \I__1146\ : Odrv4
    port map (
            O => \N__5123\,
            I => \led_blink_inst.r_Count_4Z0Z_1\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5120\,
            I => \led_blink_inst.r_Count_4Z0Z_1\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__5113\,
            I => \led_blink_inst.o_LED_43_17_cascade_\
        );

    \I__1143\ : IoInMux
    port map (
            O => \N__5110\,
            I => \N__5106\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5103\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5106\,
            I => \o_LED_4_c\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5103\,
            I => \o_LED_4_c\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5098\,
            I => \N__5095\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5095\,
            I => \led_blink_inst.r_Count_4_RNO_0Z0Z_20\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__5092\,
            I => \N__5083\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__5091\,
            I => \N__5080\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5073\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5089\,
            I => \N__5073\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5062\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5062\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5062\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5083\,
            I => \N__5062\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5080\,
            I => \N__5062\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5079\,
            I => \N__5057\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5057\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5073\,
            I => \N__5054\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5062\,
            I => \led_blink_inst.o_LED_43_17\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5057\,
            I => \led_blink_inst.o_LED_43_17\
        );

    \I__1123\ : Odrv4
    port map (
            O => \N__5054\,
            I => \led_blink_inst.o_LED_43_17\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5041\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5046\,
            I => \N__5041\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__5041\,
            I => \N__5031\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5022\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5022\
        );

    \I__1117\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5022\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5022\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5036\,
            I => \N__5015\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5035\,
            I => \N__5015\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5034\,
            I => \N__5015\
        );

    \I__1112\ : Odrv4
    port map (
            O => \N__5031\,
            I => \led_blink_inst.o_LED_43_16\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__5022\,
            I => \led_blink_inst.o_LED_43_16\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5015\,
            I => \led_blink_inst.o_LED_43_16\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__5008\,
            I => \N__5005\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5005\,
            I => \N__5002\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__5002\,
            I => \led_blink_inst.r_Count_4_RNO_0Z0Z_17\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__4999\,
            I => \N__4995\
        );

    \I__1105\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4984\
        );

    \I__1104\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4984\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__4994\,
            I => \N__4979\
        );

    \I__1102\ : InMux
    port map (
            O => \N__4993\,
            I => \N__4968\
        );

    \I__1101\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4968\
        );

    \I__1100\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4968\
        );

    \I__1099\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4968\
        );

    \I__1098\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4968\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__4984\,
            I => \N__4965\
        );

    \I__1096\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4958\
        );

    \I__1095\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4958\
        );

    \I__1094\ : InMux
    port map (
            O => \N__4979\,
            I => \N__4958\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__4968\,
            I => \led_blink_inst.o_LED_43_21\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__4965\,
            I => \led_blink_inst.o_LED_43_21\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__4958\,
            I => \led_blink_inst.o_LED_43_21\
        );

    \I__1090\ : ClkMux
    port map (
            O => \N__4951\,
            I => \N__4876\
        );

    \I__1089\ : ClkMux
    port map (
            O => \N__4950\,
            I => \N__4876\
        );

    \I__1088\ : ClkMux
    port map (
            O => \N__4949\,
            I => \N__4876\
        );

    \I__1087\ : ClkMux
    port map (
            O => \N__4948\,
            I => \N__4876\
        );

    \I__1086\ : ClkMux
    port map (
            O => \N__4947\,
            I => \N__4876\
        );

    \I__1085\ : ClkMux
    port map (
            O => \N__4946\,
            I => \N__4876\
        );

    \I__1084\ : ClkMux
    port map (
            O => \N__4945\,
            I => \N__4876\
        );

    \I__1083\ : ClkMux
    port map (
            O => \N__4944\,
            I => \N__4876\
        );

    \I__1082\ : ClkMux
    port map (
            O => \N__4943\,
            I => \N__4876\
        );

    \I__1081\ : ClkMux
    port map (
            O => \N__4942\,
            I => \N__4876\
        );

    \I__1080\ : ClkMux
    port map (
            O => \N__4941\,
            I => \N__4876\
        );

    \I__1079\ : ClkMux
    port map (
            O => \N__4940\,
            I => \N__4876\
        );

    \I__1078\ : ClkMux
    port map (
            O => \N__4939\,
            I => \N__4876\
        );

    \I__1077\ : ClkMux
    port map (
            O => \N__4938\,
            I => \N__4876\
        );

    \I__1076\ : ClkMux
    port map (
            O => \N__4937\,
            I => \N__4876\
        );

    \I__1075\ : ClkMux
    port map (
            O => \N__4936\,
            I => \N__4876\
        );

    \I__1074\ : ClkMux
    port map (
            O => \N__4935\,
            I => \N__4876\
        );

    \I__1073\ : ClkMux
    port map (
            O => \N__4934\,
            I => \N__4876\
        );

    \I__1072\ : ClkMux
    port map (
            O => \N__4933\,
            I => \N__4876\
        );

    \I__1071\ : ClkMux
    port map (
            O => \N__4932\,
            I => \N__4876\
        );

    \I__1070\ : ClkMux
    port map (
            O => \N__4931\,
            I => \N__4876\
        );

    \I__1069\ : ClkMux
    port map (
            O => \N__4930\,
            I => \N__4876\
        );

    \I__1068\ : ClkMux
    port map (
            O => \N__4929\,
            I => \N__4876\
        );

    \I__1067\ : ClkMux
    port map (
            O => \N__4928\,
            I => \N__4876\
        );

    \I__1066\ : ClkMux
    port map (
            O => \N__4927\,
            I => \N__4876\
        );

    \I__1065\ : GlobalMux
    port map (
            O => \N__4876\,
            I => \N__4873\
        );

    \I__1064\ : gio2CtrlBuf
    port map (
            O => \N__4873\,
            I => \i_Clk_c_g\
        );

    \I__1063\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4866\
        );

    \I__1062\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4863\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__4866\,
            I => \N__4860\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__4863\,
            I => \led_blink_inst.r_Count_4Z0Z_12\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__4860\,
            I => \led_blink_inst.r_Count_4Z0Z_12\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__4855\,
            I => \N__4851\
        );

    \I__1057\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4848\
        );

    \I__1056\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4845\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__4848\,
            I => \led_blink_inst.r_Count_4Z0Z_16\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__4845\,
            I => \led_blink_inst.r_Count_4Z0Z_16\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__4840\,
            I => \N__4836\
        );

    \I__1052\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4833\
        );

    \I__1051\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4830\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__4833\,
            I => \led_blink_inst.r_Count_4Z0Z_17\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__4830\,
            I => \led_blink_inst.r_Count_4Z0Z_17\
        );

    \I__1048\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4821\
        );

    \I__1047\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4818\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__4821\,
            I => \led_blink_inst.r_Count_4Z0Z_20\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__4818\,
            I => \led_blink_inst.r_Count_4Z0Z_20\
        );

    \I__1044\ : InMux
    port map (
            O => \N__4813\,
            I => \N__4810\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__4810\,
            I => \led_blink_inst.o_LED_43_15\
        );

    \I__1042\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4804\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__4804\,
            I => \led_blink_inst.r_Count_4_RNO_0Z0Z_9\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4797\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4794\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__4797\,
            I => \led_blink_inst.r_Count_4Z0Z_6\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__4794\,
            I => \led_blink_inst.r_Count_4Z0Z_6\
        );

    \I__1036\ : InMux
    port map (
            O => \N__4789\,
            I => \N__4785\
        );

    \I__1035\ : InMux
    port map (
            O => \N__4788\,
            I => \N__4782\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__4785\,
            I => \led_blink_inst.r_Count_4Z0Z_9\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__4782\,
            I => \led_blink_inst.r_Count_4Z0Z_9\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__4777\,
            I => \N__4774\
        );

    \I__1031\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4770\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4767\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__4770\,
            I => \led_blink_inst.r_Count_4Z0Z_7\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4767\,
            I => \led_blink_inst.r_Count_4Z0Z_7\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4758\
        );

    \I__1026\ : InMux
    port map (
            O => \N__4761\,
            I => \N__4755\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__4758\,
            I => \led_blink_inst.r_Count_4Z0Z_4\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__4755\,
            I => \led_blink_inst.r_Count_4Z0Z_4\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__4750\,
            I => \N__4746\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4743\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4740\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__4743\,
            I => \led_blink_inst.r_Count_4Z0Z_8\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__4740\,
            I => \led_blink_inst.r_Count_4Z0Z_8\
        );

    \I__1018\ : InMux
    port map (
            O => \N__4735\,
            I => \N__4731\
        );

    \I__1017\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4728\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__4731\,
            I => \led_blink_inst.r_Count_4Z0Z_10\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__4728\,
            I => \led_blink_inst.r_Count_4Z0Z_10\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__4723\,
            I => \N__4719\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__4722\,
            I => \N__4716\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4713\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4710\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4713\,
            I => \led_blink_inst.r_Count_4Z0Z_13\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__4710\,
            I => \led_blink_inst.r_Count_4Z0Z_13\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__4705\,
            I => \N__4701\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4704\,
            I => \N__4698\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4701\,
            I => \N__4695\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4698\,
            I => \led_blink_inst.r_Count_4Z0Z_5\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4695\,
            I => \led_blink_inst.r_Count_4Z0Z_5\
        );

    \I__1003\ : CascadeMux
    port map (
            O => \N__4690\,
            I => \led_blink_inst.o_LED_43_16_cascade_\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4684\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__4684\,
            I => \led_blink_inst.r_Count_4_RNO_0Z0Z_16\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__4681\,
            I => \N__4678\
        );

    \I__999\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4675\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4675\,
            I => \led_blink_inst.r_Count_4_RNO_0Z0Z_12\
        );

    \I__997\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4669\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__4669\,
            I => \N__4665\
        );

    \I__995\ : InMux
    port map (
            O => \N__4668\,
            I => \N__4662\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__4665\,
            I => \led_blink_inst.r_Count_4Z0Z_14\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4662\,
            I => \led_blink_inst.r_Count_4Z0Z_14\
        );

    \I__992\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4653\
        );

    \I__991\ : InMux
    port map (
            O => \N__4656\,
            I => \N__4650\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4653\,
            I => \led_blink_inst.r_Count_4Z0Z_23\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4650\,
            I => \led_blink_inst.r_Count_4Z0Z_23\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__4645\,
            I => \N__4641\
        );

    \I__987\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4638\
        );

    \I__986\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4635\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4638\,
            I => \led_blink_inst.r_Count_4Z0Z_21\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4635\,
            I => \led_blink_inst.r_Count_4Z0Z_21\
        );

    \I__983\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4626\
        );

    \I__982\ : InMux
    port map (
            O => \N__4629\,
            I => \N__4623\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4626\,
            I => \led_blink_inst.r_Count_4Z0Z_3\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4623\,
            I => \led_blink_inst.r_Count_4Z0Z_3\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__4618\,
            I => \N__4614\
        );

    \I__978\ : InMux
    port map (
            O => \N__4617\,
            I => \N__4611\
        );

    \I__977\ : InMux
    port map (
            O => \N__4614\,
            I => \N__4608\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4611\,
            I => \led_blink_inst.r_Count_3Z0Z_18\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__4608\,
            I => \led_blink_inst.r_Count_3Z0Z_18\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__4603\,
            I => \N__4600\
        );

    \I__973\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4597\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4597\,
            I => \led_blink_inst.r_Count_3_RNO_0Z0Z_18\
        );

    \I__971\ : InMux
    port map (
            O => \N__4594\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_17\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__4591\,
            I => \N__4587\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__4590\,
            I => \N__4584\
        );

    \I__968\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4581\
        );

    \I__967\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4578\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4581\,
            I => \led_blink_inst.r_Count_3Z0Z_19\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__4578\,
            I => \led_blink_inst.r_Count_3Z0Z_19\
        );

    \I__964\ : InMux
    port map (
            O => \N__4573\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_18\
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__4570\,
            I => \N__4566\
        );

    \I__962\ : InMux
    port map (
            O => \N__4569\,
            I => \N__4563\
        );

    \I__961\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4560\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4563\,
            I => \led_blink_inst.r_Count_3Z0Z_20\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4560\,
            I => \led_blink_inst.r_Count_3Z0Z_20\
        );

    \I__958\ : InMux
    port map (
            O => \N__4555\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_19\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__4552\,
            I => \N__4548\
        );

    \I__956\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4545\
        );

    \I__955\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4542\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4545\,
            I => \led_blink_inst.r_Count_3Z0Z_21\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4542\,
            I => \led_blink_inst.r_Count_3Z0Z_21\
        );

    \I__952\ : InMux
    port map (
            O => \N__4537\,
            I => \N__4534\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4534\,
            I => \led_blink_inst.r_Count_3_RNO_0Z0Z_21\
        );

    \I__950\ : InMux
    port map (
            O => \N__4531\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_20\
        );

    \I__949\ : CascadeMux
    port map (
            O => \N__4528\,
            I => \N__4524\
        );

    \I__948\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4521\
        );

    \I__947\ : InMux
    port map (
            O => \N__4524\,
            I => \N__4518\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4521\,
            I => \led_blink_inst.r_Count_3Z0Z_22\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4518\,
            I => \led_blink_inst.r_Count_3Z0Z_22\
        );

    \I__944\ : InMux
    port map (
            O => \N__4513\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_21\
        );

    \I__943\ : InMux
    port map (
            O => \N__4510\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_22\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__4507\,
            I => \N__4504\
        );

    \I__941\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4500\
        );

    \I__940\ : InMux
    port map (
            O => \N__4503\,
            I => \N__4497\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4500\,
            I => \N__4494\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4497\,
            I => \led_blink_inst.r_Count_3Z0Z_23\
        );

    \I__937\ : Odrv4
    port map (
            O => \N__4494\,
            I => \led_blink_inst.r_Count_3Z0Z_23\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__4489\,
            I => \N__4486\
        );

    \I__935\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4483\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4483\,
            I => \N__4480\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__4480\,
            I => \led_blink_inst.r_Count_4_RNO_0Z0Z_4\
        );

    \I__932\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4474\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4474\,
            I => \led_blink_inst.r_Count_4_RNO_0Z0Z_7\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__4471\,
            I => \N__4468\
        );

    \I__929\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4465\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4465\,
            I => \led_blink_inst.r_Count_4_RNO_0Z0Z_6\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__4462\,
            I => \N__4458\
        );

    \I__926\ : CascadeMux
    port map (
            O => \N__4461\,
            I => \N__4455\
        );

    \I__925\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4452\
        );

    \I__924\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4449\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4452\,
            I => \led_blink_inst.r_Count_3Z0Z_10\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4449\,
            I => \led_blink_inst.r_Count_3Z0Z_10\
        );

    \I__921\ : InMux
    port map (
            O => \N__4444\,
            I => \N__4441\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4441\,
            I => \led_blink_inst.r_Count_3_RNO_0Z0Z_10\
        );

    \I__919\ : InMux
    port map (
            O => \N__4438\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_9\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__4435\,
            I => \N__4431\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__4434\,
            I => \N__4428\
        );

    \I__916\ : InMux
    port map (
            O => \N__4431\,
            I => \N__4425\
        );

    \I__915\ : InMux
    port map (
            O => \N__4428\,
            I => \N__4422\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4425\,
            I => \led_blink_inst.r_Count_3Z0Z_11\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4422\,
            I => \led_blink_inst.r_Count_3Z0Z_11\
        );

    \I__912\ : InMux
    port map (
            O => \N__4417\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_10\
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__4414\,
            I => \N__4410\
        );

    \I__910\ : InMux
    port map (
            O => \N__4413\,
            I => \N__4407\
        );

    \I__909\ : InMux
    port map (
            O => \N__4410\,
            I => \N__4404\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4407\,
            I => \led_blink_inst.r_Count_3Z0Z_12\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4404\,
            I => \led_blink_inst.r_Count_3Z0Z_12\
        );

    \I__906\ : InMux
    port map (
            O => \N__4399\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_11\
        );

    \I__905\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4392\
        );

    \I__904\ : InMux
    port map (
            O => \N__4395\,
            I => \N__4389\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4392\,
            I => \led_blink_inst.r_Count_3Z0Z_13\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4389\,
            I => \led_blink_inst.r_Count_3Z0Z_13\
        );

    \I__901\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4381\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4381\,
            I => \led_blink_inst.r_Count_3_RNO_0Z0Z_13\
        );

    \I__899\ : InMux
    port map (
            O => \N__4378\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_12\
        );

    \I__898\ : InMux
    port map (
            O => \N__4375\,
            I => \N__4372\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4372\,
            I => \N__4368\
        );

    \I__896\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4365\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__4368\,
            I => \led_blink_inst.r_Count_3Z0Z_14\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4365\,
            I => \led_blink_inst.r_Count_3Z0Z_14\
        );

    \I__893\ : InMux
    port map (
            O => \N__4360\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_13\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__4357\,
            I => \N__4353\
        );

    \I__891\ : InMux
    port map (
            O => \N__4356\,
            I => \N__4350\
        );

    \I__890\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4347\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4350\,
            I => \led_blink_inst.r_Count_3Z0Z_15\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4347\,
            I => \led_blink_inst.r_Count_3Z0Z_15\
        );

    \I__887\ : InMux
    port map (
            O => \N__4342\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_14\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__4339\,
            I => \N__4335\
        );

    \I__885\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4332\
        );

    \I__884\ : InMux
    port map (
            O => \N__4335\,
            I => \N__4329\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4332\,
            I => \led_blink_inst.r_Count_3Z0Z_16\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4329\,
            I => \led_blink_inst.r_Count_3Z0Z_16\
        );

    \I__881\ : InMux
    port map (
            O => \N__4324\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_15\
        );

    \I__880\ : InMux
    port map (
            O => \N__4321\,
            I => \N__4317\
        );

    \I__879\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4314\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4317\,
            I => \led_blink_inst.r_Count_3Z0Z_17\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4314\,
            I => \led_blink_inst.r_Count_3Z0Z_17\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__4309\,
            I => \N__4306\
        );

    \I__875\ : InMux
    port map (
            O => \N__4306\,
            I => \N__4303\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4303\,
            I => \led_blink_inst.r_Count_3_RNO_0Z0Z_17\
        );

    \I__873\ : InMux
    port map (
            O => \N__4300\,
            I => \bfn_12_5_0_\
        );

    \I__872\ : InMux
    port map (
            O => \N__4297\,
            I => \N__4293\
        );

    \I__871\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4290\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4293\,
            I => \led_blink_inst.r_Count_3Z0Z_2\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4290\,
            I => \led_blink_inst.r_Count_3Z0Z_2\
        );

    \I__868\ : InMux
    port map (
            O => \N__4285\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_1\
        );

    \I__867\ : InMux
    port map (
            O => \N__4282\,
            I => \N__4278\
        );

    \I__866\ : InMux
    port map (
            O => \N__4281\,
            I => \N__4275\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4278\,
            I => \led_blink_inst.r_Count_3Z0Z_3\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4275\,
            I => \led_blink_inst.r_Count_3Z0Z_3\
        );

    \I__863\ : InMux
    port map (
            O => \N__4270\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_2\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__4267\,
            I => \N__4263\
        );

    \I__861\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4260\
        );

    \I__860\ : InMux
    port map (
            O => \N__4263\,
            I => \N__4257\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4260\,
            I => \led_blink_inst.r_Count_3Z0Z_4\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4257\,
            I => \led_blink_inst.r_Count_3Z0Z_4\
        );

    \I__857\ : InMux
    port map (
            O => \N__4252\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_3\
        );

    \I__856\ : InMux
    port map (
            O => \N__4249\,
            I => \N__4245\
        );

    \I__855\ : InMux
    port map (
            O => \N__4248\,
            I => \N__4242\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4245\,
            I => \led_blink_inst.r_Count_3Z0Z_5\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4242\,
            I => \led_blink_inst.r_Count_3Z0Z_5\
        );

    \I__852\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4234\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4234\,
            I => \led_blink_inst.r_Count_3_RNO_0Z0Z_5\
        );

    \I__850\ : InMux
    port map (
            O => \N__4231\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_4\
        );

    \I__849\ : InMux
    port map (
            O => \N__4228\,
            I => \N__4225\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4225\,
            I => \N__4221\
        );

    \I__847\ : InMux
    port map (
            O => \N__4224\,
            I => \N__4218\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__4221\,
            I => \led_blink_inst.r_Count_3Z0Z_6\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4218\,
            I => \led_blink_inst.r_Count_3Z0Z_6\
        );

    \I__844\ : InMux
    port map (
            O => \N__4213\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_5\
        );

    \I__843\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4207\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4207\,
            I => \N__4203\
        );

    \I__841\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4200\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__4203\,
            I => \led_blink_inst.r_Count_3Z0Z_7\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4200\,
            I => \led_blink_inst.r_Count_3Z0Z_7\
        );

    \I__838\ : InMux
    port map (
            O => \N__4195\,
            I => \N__4192\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4192\,
            I => \led_blink_inst.r_Count_3_RNO_0Z0Z_7\
        );

    \I__836\ : InMux
    port map (
            O => \N__4189\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_6\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__4186\,
            I => \N__4182\
        );

    \I__834\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4179\
        );

    \I__833\ : InMux
    port map (
            O => \N__4182\,
            I => \N__4176\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4179\,
            I => \led_blink_inst.r_Count_3Z0Z_8\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4176\,
            I => \led_blink_inst.r_Count_3Z0Z_8\
        );

    \I__830\ : CascadeMux
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__829\ : InMux
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4165\,
            I => \N__4162\
        );

    \I__827\ : Odrv4
    port map (
            O => \N__4162\,
            I => \led_blink_inst.r_Count_3_RNO_0Z0Z_8\
        );

    \I__826\ : InMux
    port map (
            O => \N__4159\,
            I => \led_blink_inst.un2_r_Count_3_1_cry_7\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__4156\,
            I => \N__4152\
        );

    \I__824\ : InMux
    port map (
            O => \N__4155\,
            I => \N__4149\
        );

    \I__823\ : InMux
    port map (
            O => \N__4152\,
            I => \N__4146\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4149\,
            I => \led_blink_inst.r_Count_3Z0Z_9\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4146\,
            I => \led_blink_inst.r_Count_3Z0Z_9\
        );

    \I__820\ : InMux
    port map (
            O => \N__4141\,
            I => \bfn_12_4_0_\
        );

    \I__819\ : InMux
    port map (
            O => \N__4138\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_15\
        );

    \I__818\ : InMux
    port map (
            O => \N__4135\,
            I => \bfn_11_8_0_\
        );

    \I__817\ : InMux
    port map (
            O => \N__4132\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_17\
        );

    \I__816\ : InMux
    port map (
            O => \N__4129\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_18\
        );

    \I__815\ : InMux
    port map (
            O => \N__4126\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_19\
        );

    \I__814\ : InMux
    port map (
            O => \N__4123\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_20\
        );

    \I__813\ : InMux
    port map (
            O => \N__4120\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_21\
        );

    \I__812\ : InMux
    port map (
            O => \N__4117\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_22\
        );

    \I__811\ : InMux
    port map (
            O => \N__4114\,
            I => \N__4107\
        );

    \I__810\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4107\
        );

    \I__809\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4104\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4107\,
            I => \led_blink_inst.r_Count_3Z0Z_1\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4104\,
            I => \led_blink_inst.r_Count_3Z0Z_1\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__4099\,
            I => \N__4093\
        );

    \I__805\ : InMux
    port map (
            O => \N__4098\,
            I => \N__4090\
        );

    \I__804\ : InMux
    port map (
            O => \N__4097\,
            I => \N__4085\
        );

    \I__803\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4085\
        );

    \I__802\ : InMux
    port map (
            O => \N__4093\,
            I => \N__4082\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4090\,
            I => \led_blink_inst.r_Count_3Z0Z_0\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4085\,
            I => \led_blink_inst.r_Count_3Z0Z_0\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4082\,
            I => \led_blink_inst.r_Count_3Z0Z_0\
        );

    \I__798\ : InMux
    port map (
            O => \N__4075\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_6\
        );

    \I__797\ : InMux
    port map (
            O => \N__4072\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_7\
        );

    \I__796\ : InMux
    port map (
            O => \N__4069\,
            I => \bfn_11_7_0_\
        );

    \I__795\ : InMux
    port map (
            O => \N__4066\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_9\
        );

    \I__794\ : InMux
    port map (
            O => \N__4063\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_10\
        );

    \I__793\ : InMux
    port map (
            O => \N__4060\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_11\
        );

    \I__792\ : InMux
    port map (
            O => \N__4057\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_12\
        );

    \I__791\ : InMux
    port map (
            O => \N__4054\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_13\
        );

    \I__790\ : InMux
    port map (
            O => \N__4051\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_14\
        );

    \I__789\ : InMux
    port map (
            O => \N__4048\,
            I => \N__4045\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4045\,
            I => \led_blink_inst.o_LED_33_15\
        );

    \I__787\ : InMux
    port map (
            O => \N__4042\,
            I => \N__4029\
        );

    \I__786\ : InMux
    port map (
            O => \N__4041\,
            I => \N__4029\
        );

    \I__785\ : InMux
    port map (
            O => \N__4040\,
            I => \N__4029\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__4039\,
            I => \N__4024\
        );

    \I__783\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4016\
        );

    \I__782\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4016\
        );

    \I__781\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4016\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4029\,
            I => \N__4013\
        );

    \I__779\ : InMux
    port map (
            O => \N__4028\,
            I => \N__4006\
        );

    \I__778\ : InMux
    port map (
            O => \N__4027\,
            I => \N__4006\
        );

    \I__777\ : InMux
    port map (
            O => \N__4024\,
            I => \N__4006\
        );

    \I__776\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4003\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4016\,
            I => \led_blink_inst.o_LED_33_17\
        );

    \I__774\ : Odrv4
    port map (
            O => \N__4013\,
            I => \led_blink_inst.o_LED_33_17\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4006\,
            I => \led_blink_inst.o_LED_33_17\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__4003\,
            I => \led_blink_inst.o_LED_33_17\
        );

    \I__771\ : InMux
    port map (
            O => \N__3994\,
            I => \N__3979\
        );

    \I__770\ : InMux
    port map (
            O => \N__3993\,
            I => \N__3979\
        );

    \I__769\ : InMux
    port map (
            O => \N__3992\,
            I => \N__3979\
        );

    \I__768\ : InMux
    port map (
            O => \N__3991\,
            I => \N__3972\
        );

    \I__767\ : InMux
    port map (
            O => \N__3990\,
            I => \N__3972\
        );

    \I__766\ : InMux
    port map (
            O => \N__3989\,
            I => \N__3972\
        );

    \I__765\ : InMux
    port map (
            O => \N__3988\,
            I => \N__3965\
        );

    \I__764\ : InMux
    port map (
            O => \N__3987\,
            I => \N__3965\
        );

    \I__763\ : InMux
    port map (
            O => \N__3986\,
            I => \N__3965\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__3979\,
            I => \led_blink_inst.o_LED_33_16\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__3972\,
            I => \led_blink_inst.o_LED_33_16\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__3965\,
            I => \led_blink_inst.o_LED_33_16\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__3958\,
            I => \N__3951\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__3957\,
            I => \N__3948\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__3956\,
            I => \N__3943\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__3955\,
            I => \N__3938\
        );

    \I__755\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3935\
        );

    \I__754\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3930\
        );

    \I__753\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3930\
        );

    \I__752\ : InMux
    port map (
            O => \N__3947\,
            I => \N__3923\
        );

    \I__751\ : InMux
    port map (
            O => \N__3946\,
            I => \N__3923\
        );

    \I__750\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3923\
        );

    \I__749\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3916\
        );

    \I__748\ : InMux
    port map (
            O => \N__3941\,
            I => \N__3916\
        );

    \I__747\ : InMux
    port map (
            O => \N__3938\,
            I => \N__3916\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__3935\,
            I => \led_blink_inst.o_LED_33_21\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3930\,
            I => \led_blink_inst.o_LED_33_21\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__3923\,
            I => \led_blink_inst.o_LED_33_21\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3916\,
            I => \led_blink_inst.o_LED_33_21\
        );

    \I__742\ : InMux
    port map (
            O => \N__3907\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_1\
        );

    \I__741\ : InMux
    port map (
            O => \N__3904\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_2\
        );

    \I__740\ : InMux
    port map (
            O => \N__3901\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_3\
        );

    \I__739\ : InMux
    port map (
            O => \N__3898\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_4\
        );

    \I__738\ : InMux
    port map (
            O => \N__3895\,
            I => \led_blink_inst.un2_r_Count_4_1_cry_5\
        );

    \I__737\ : InMux
    port map (
            O => \N__3892\,
            I => \N__3889\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3889\,
            I => \N__3886\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__3886\,
            I => \led_blink_inst.o_LED_33_14\
        );

    \I__734\ : InMux
    port map (
            O => \N__3883\,
            I => \N__3880\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3880\,
            I => \led_blink_inst.o_LED_33_13\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__3877\,
            I => \led_blink_inst.o_LED_33_12_cascade_\
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__3874\,
            I => \led_blink_inst.o_LED_33_21_cascade_\
        );

    \I__730\ : IoInMux
    port map (
            O => \N__3871\,
            I => \N__3868\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3868\,
            I => \N__3864\
        );

    \I__728\ : InMux
    port map (
            O => \N__3867\,
            I => \N__3861\
        );

    \I__727\ : Span4Mux_s1_h
    port map (
            O => \N__3864\,
            I => \N__3858\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__3861\,
            I => \N__3855\
        );

    \I__725\ : Odrv4
    port map (
            O => \N__3858\,
            I => \o_LED_3_c\
        );

    \I__724\ : Odrv4
    port map (
            O => \N__3855\,
            I => \o_LED_3_c\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__3850\,
            I => \led_blink_inst.o_LED_33_16_cascade_\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__3847\,
            I => \N__3844\
        );

    \I__721\ : InMux
    port map (
            O => \N__3844\,
            I => \N__3840\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__3843\,
            I => \N__3837\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3840\,
            I => \N__3834\
        );

    \I__718\ : InMux
    port map (
            O => \N__3837\,
            I => \N__3831\
        );

    \I__717\ : Odrv4
    port map (
            O => \N__3834\,
            I => \led_blink_inst.r_Count_2Z0Z_21\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3831\,
            I => \led_blink_inst.r_Count_2Z0Z_21\
        );

    \I__715\ : InMux
    port map (
            O => \N__3826\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_20\
        );

    \I__714\ : InMux
    port map (
            O => \N__3823\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_21\
        );

    \I__713\ : InMux
    port map (
            O => \N__3820\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_22\
        );

    \I__712\ : InMux
    port map (
            O => \N__3817\,
            I => \N__3813\
        );

    \I__711\ : InMux
    port map (
            O => \N__3816\,
            I => \N__3810\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3813\,
            I => \N__3807\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3810\,
            I => \led_blink_inst.r_Count_2Z0Z_23\
        );

    \I__708\ : Odrv12
    port map (
            O => \N__3807\,
            I => \led_blink_inst.r_Count_2Z0Z_23\
        );

    \I__707\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3798\
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__3801\,
            I => \N__3783\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3798\,
            I => \N__3780\
        );

    \I__704\ : InMux
    port map (
            O => \N__3797\,
            I => \N__3767\
        );

    \I__703\ : InMux
    port map (
            O => \N__3796\,
            I => \N__3767\
        );

    \I__702\ : InMux
    port map (
            O => \N__3795\,
            I => \N__3767\
        );

    \I__701\ : InMux
    port map (
            O => \N__3794\,
            I => \N__3767\
        );

    \I__700\ : InMux
    port map (
            O => \N__3793\,
            I => \N__3767\
        );

    \I__699\ : InMux
    port map (
            O => \N__3792\,
            I => \N__3767\
        );

    \I__698\ : InMux
    port map (
            O => \N__3791\,
            I => \N__3764\
        );

    \I__697\ : InMux
    port map (
            O => \N__3790\,
            I => \N__3757\
        );

    \I__696\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3757\
        );

    \I__695\ : InMux
    port map (
            O => \N__3788\,
            I => \N__3757\
        );

    \I__694\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3750\
        );

    \I__693\ : InMux
    port map (
            O => \N__3786\,
            I => \N__3750\
        );

    \I__692\ : InMux
    port map (
            O => \N__3783\,
            I => \N__3750\
        );

    \I__691\ : Odrv12
    port map (
            O => \N__3780\,
            I => \led_blink_inst.o_LED_23_17\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3767\,
            I => \led_blink_inst.o_LED_23_17\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3764\,
            I => \led_blink_inst.o_LED_23_17\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3757\,
            I => \led_blink_inst.o_LED_23_17\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3750\,
            I => \led_blink_inst.o_LED_23_17\
        );

    \I__686\ : InMux
    port map (
            O => \N__3739\,
            I => \N__3736\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__684\ : Span4Mux_v
    port map (
            O => \N__3733\,
            I => \N__3718\
        );

    \I__683\ : InMux
    port map (
            O => \N__3732\,
            I => \N__3705\
        );

    \I__682\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3705\
        );

    \I__681\ : InMux
    port map (
            O => \N__3730\,
            I => \N__3705\
        );

    \I__680\ : InMux
    port map (
            O => \N__3729\,
            I => \N__3705\
        );

    \I__679\ : InMux
    port map (
            O => \N__3728\,
            I => \N__3705\
        );

    \I__678\ : InMux
    port map (
            O => \N__3727\,
            I => \N__3705\
        );

    \I__677\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3698\
        );

    \I__676\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3698\
        );

    \I__675\ : InMux
    port map (
            O => \N__3724\,
            I => \N__3698\
        );

    \I__674\ : InMux
    port map (
            O => \N__3723\,
            I => \N__3691\
        );

    \I__673\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3691\
        );

    \I__672\ : InMux
    port map (
            O => \N__3721\,
            I => \N__3691\
        );

    \I__671\ : Odrv4
    port map (
            O => \N__3718\,
            I => \led_blink_inst.o_LED_23_16\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3705\,
            I => \led_blink_inst.o_LED_23_16\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3698\,
            I => \led_blink_inst.o_LED_23_16\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3691\,
            I => \led_blink_inst.o_LED_23_16\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__3682\,
            I => \N__3679\
        );

    \I__666\ : InMux
    port map (
            O => \N__3679\,
            I => \N__3676\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3676\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_22\
        );

    \I__664\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3666\
        );

    \I__663\ : CascadeMux
    port map (
            O => \N__3672\,
            I => \N__3661\
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__3671\,
            I => \N__3657\
        );

    \I__661\ : CascadeMux
    port map (
            O => \N__3670\,
            I => \N__3652\
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__3669\,
            I => \N__3647\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3666\,
            I => \N__3643\
        );

    \I__658\ : InMux
    port map (
            O => \N__3665\,
            I => \N__3630\
        );

    \I__657\ : InMux
    port map (
            O => \N__3664\,
            I => \N__3630\
        );

    \I__656\ : InMux
    port map (
            O => \N__3661\,
            I => \N__3630\
        );

    \I__655\ : InMux
    port map (
            O => \N__3660\,
            I => \N__3630\
        );

    \I__654\ : InMux
    port map (
            O => \N__3657\,
            I => \N__3630\
        );

    \I__653\ : InMux
    port map (
            O => \N__3656\,
            I => \N__3630\
        );

    \I__652\ : InMux
    port map (
            O => \N__3655\,
            I => \N__3627\
        );

    \I__651\ : InMux
    port map (
            O => \N__3652\,
            I => \N__3620\
        );

    \I__650\ : InMux
    port map (
            O => \N__3651\,
            I => \N__3620\
        );

    \I__649\ : InMux
    port map (
            O => \N__3650\,
            I => \N__3620\
        );

    \I__648\ : InMux
    port map (
            O => \N__3647\,
            I => \N__3615\
        );

    \I__647\ : InMux
    port map (
            O => \N__3646\,
            I => \N__3615\
        );

    \I__646\ : Odrv4
    port map (
            O => \N__3643\,
            I => \led_blink_inst.o_LED_23_21\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3630\,
            I => \led_blink_inst.o_LED_23_21\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3627\,
            I => \led_blink_inst.o_LED_23_21\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3620\,
            I => \led_blink_inst.o_LED_23_21\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3615\,
            I => \led_blink_inst.o_LED_23_21\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__3604\,
            I => \N__3601\
        );

    \I__640\ : InMux
    port map (
            O => \N__3601\,
            I => \N__3598\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__3598\,
            I => \N__3595\
        );

    \I__638\ : Span4Mux_h
    port map (
            O => \N__3595\,
            I => \N__3591\
        );

    \I__637\ : InMux
    port map (
            O => \N__3594\,
            I => \N__3588\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__3591\,
            I => \led_blink_inst.r_Count_2Z0Z_22\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3588\,
            I => \led_blink_inst.r_Count_2Z0Z_22\
        );

    \I__634\ : CascadeMux
    port map (
            O => \N__3583\,
            I => \N__3580\
        );

    \I__633\ : InMux
    port map (
            O => \N__3580\,
            I => \N__3577\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3577\,
            I => \N__3573\
        );

    \I__631\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3570\
        );

    \I__630\ : Odrv12
    port map (
            O => \N__3573\,
            I => \led_blink_inst.r_Count_2Z0Z_13\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3570\,
            I => \led_blink_inst.r_Count_2Z0Z_13\
        );

    \I__628\ : InMux
    port map (
            O => \N__3565\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_12\
        );

    \I__627\ : InMux
    port map (
            O => \N__3562\,
            I => \N__3558\
        );

    \I__626\ : InMux
    port map (
            O => \N__3561\,
            I => \N__3555\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3558\,
            I => \led_blink_inst.r_Count_2Z0Z_14\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3555\,
            I => \led_blink_inst.r_Count_2Z0Z_14\
        );

    \I__623\ : InMux
    port map (
            O => \N__3550\,
            I => \N__3547\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3547\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_14\
        );

    \I__621\ : InMux
    port map (
            O => \N__3544\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_13\
        );

    \I__620\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3537\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__3540\,
            I => \N__3534\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3537\,
            I => \N__3531\
        );

    \I__617\ : InMux
    port map (
            O => \N__3534\,
            I => \N__3528\
        );

    \I__616\ : Odrv4
    port map (
            O => \N__3531\,
            I => \led_blink_inst.r_Count_2Z0Z_15\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3528\,
            I => \led_blink_inst.r_Count_2Z0Z_15\
        );

    \I__614\ : InMux
    port map (
            O => \N__3523\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_14\
        );

    \I__613\ : InMux
    port map (
            O => \N__3520\,
            I => \N__3516\
        );

    \I__612\ : InMux
    port map (
            O => \N__3519\,
            I => \N__3513\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3516\,
            I => \N__3510\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3513\,
            I => \led_blink_inst.r_Count_2Z0Z_16\
        );

    \I__609\ : Odrv12
    port map (
            O => \N__3510\,
            I => \led_blink_inst.r_Count_2Z0Z_16\
        );

    \I__608\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3502\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3502\,
            I => \N__3499\
        );

    \I__606\ : Odrv12
    port map (
            O => \N__3499\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_16\
        );

    \I__605\ : InMux
    port map (
            O => \N__3496\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_15\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__3493\,
            I => \N__3490\
        );

    \I__603\ : InMux
    port map (
            O => \N__3490\,
            I => \N__3486\
        );

    \I__602\ : InMux
    port map (
            O => \N__3489\,
            I => \N__3483\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3486\,
            I => \N__3480\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3483\,
            I => \led_blink_inst.r_Count_2Z0Z_17\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__3480\,
            I => \led_blink_inst.r_Count_2Z0Z_17\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__3475\,
            I => \N__3472\
        );

    \I__597\ : InMux
    port map (
            O => \N__3472\,
            I => \N__3469\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3469\,
            I => \N__3466\
        );

    \I__595\ : Span4Mux_h
    port map (
            O => \N__3466\,
            I => \N__3463\
        );

    \I__594\ : Odrv4
    port map (
            O => \N__3463\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_17\
        );

    \I__593\ : InMux
    port map (
            O => \N__3460\,
            I => \bfn_9_8_0_\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__3457\,
            I => \N__3454\
        );

    \I__591\ : InMux
    port map (
            O => \N__3454\,
            I => \N__3450\
        );

    \I__590\ : InMux
    port map (
            O => \N__3453\,
            I => \N__3447\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3450\,
            I => \N__3444\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3447\,
            I => \led_blink_inst.r_Count_2Z0Z_18\
        );

    \I__587\ : Odrv4
    port map (
            O => \N__3444\,
            I => \led_blink_inst.r_Count_2Z0Z_18\
        );

    \I__586\ : InMux
    port map (
            O => \N__3439\,
            I => \N__3436\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3436\,
            I => \N__3433\
        );

    \I__584\ : Odrv4
    port map (
            O => \N__3433\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_18\
        );

    \I__583\ : InMux
    port map (
            O => \N__3430\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_17\
        );

    \I__582\ : InMux
    port map (
            O => \N__3427\,
            I => \N__3423\
        );

    \I__581\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3420\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3423\,
            I => \N__3417\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3420\,
            I => \led_blink_inst.r_Count_2Z0Z_19\
        );

    \I__578\ : Odrv4
    port map (
            O => \N__3417\,
            I => \led_blink_inst.r_Count_2Z0Z_19\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__3412\,
            I => \N__3409\
        );

    \I__576\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3406\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3406\,
            I => \N__3403\
        );

    \I__574\ : Odrv4
    port map (
            O => \N__3403\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_19\
        );

    \I__573\ : InMux
    port map (
            O => \N__3400\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_18\
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__3397\,
            I => \N__3394\
        );

    \I__571\ : InMux
    port map (
            O => \N__3394\,
            I => \N__3390\
        );

    \I__570\ : InMux
    port map (
            O => \N__3393\,
            I => \N__3387\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3390\,
            I => \N__3384\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3387\,
            I => \led_blink_inst.r_Count_2Z0Z_20\
        );

    \I__567\ : Odrv4
    port map (
            O => \N__3384\,
            I => \led_blink_inst.r_Count_2Z0Z_20\
        );

    \I__566\ : CascadeMux
    port map (
            O => \N__3379\,
            I => \N__3376\
        );

    \I__565\ : InMux
    port map (
            O => \N__3376\,
            I => \N__3373\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__3373\,
            I => \N__3370\
        );

    \I__563\ : Odrv4
    port map (
            O => \N__3370\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_20\
        );

    \I__562\ : InMux
    port map (
            O => \N__3367\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_19\
        );

    \I__561\ : InMux
    port map (
            O => \N__3364\,
            I => \N__3360\
        );

    \I__560\ : InMux
    port map (
            O => \N__3363\,
            I => \N__3357\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3360\,
            I => \led_blink_inst.r_Count_2Z0Z_5\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3357\,
            I => \led_blink_inst.r_Count_2Z0Z_5\
        );

    \I__557\ : InMux
    port map (
            O => \N__3352\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_4\
        );

    \I__556\ : InMux
    port map (
            O => \N__3349\,
            I => \N__3345\
        );

    \I__555\ : InMux
    port map (
            O => \N__3348\,
            I => \N__3342\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3345\,
            I => \led_blink_inst.r_Count_2Z0Z_6\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3342\,
            I => \led_blink_inst.r_Count_2Z0Z_6\
        );

    \I__552\ : InMux
    port map (
            O => \N__3337\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_5\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__3334\,
            I => \N__3330\
        );

    \I__550\ : InMux
    port map (
            O => \N__3333\,
            I => \N__3327\
        );

    \I__549\ : InMux
    port map (
            O => \N__3330\,
            I => \N__3324\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3327\,
            I => \led_blink_inst.r_Count_2Z0Z_7\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3324\,
            I => \led_blink_inst.r_Count_2Z0Z_7\
        );

    \I__546\ : InMux
    port map (
            O => \N__3319\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_6\
        );

    \I__545\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3312\
        );

    \I__544\ : InMux
    port map (
            O => \N__3315\,
            I => \N__3309\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3312\,
            I => \led_blink_inst.r_Count_2Z0Z_8\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3309\,
            I => \led_blink_inst.r_Count_2Z0Z_8\
        );

    \I__541\ : InMux
    port map (
            O => \N__3304\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_7\
        );

    \I__540\ : InMux
    port map (
            O => \N__3301\,
            I => \N__3297\
        );

    \I__539\ : InMux
    port map (
            O => \N__3300\,
            I => \N__3294\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3297\,
            I => \N__3291\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3294\,
            I => \N__3288\
        );

    \I__536\ : Odrv4
    port map (
            O => \N__3291\,
            I => \led_blink_inst.r_Count_2Z0Z_9\
        );

    \I__535\ : Odrv4
    port map (
            O => \N__3288\,
            I => \led_blink_inst.r_Count_2Z0Z_9\
        );

    \I__534\ : InMux
    port map (
            O => \N__3283\,
            I => \N__3280\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3280\,
            I => \N__3277\
        );

    \I__532\ : Odrv4
    port map (
            O => \N__3277\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_9\
        );

    \I__531\ : InMux
    port map (
            O => \N__3274\,
            I => \bfn_9_7_0_\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__3271\,
            I => \N__3267\
        );

    \I__529\ : InMux
    port map (
            O => \N__3270\,
            I => \N__3264\
        );

    \I__528\ : InMux
    port map (
            O => \N__3267\,
            I => \N__3261\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3264\,
            I => \led_blink_inst.r_Count_2Z0Z_10\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3261\,
            I => \led_blink_inst.r_Count_2Z0Z_10\
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__3256\,
            I => \N__3253\
        );

    \I__524\ : InMux
    port map (
            O => \N__3253\,
            I => \N__3250\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3250\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_10\
        );

    \I__522\ : InMux
    port map (
            O => \N__3247\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_9\
        );

    \I__521\ : CascadeMux
    port map (
            O => \N__3244\,
            I => \N__3240\
        );

    \I__520\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3237\
        );

    \I__519\ : InMux
    port map (
            O => \N__3240\,
            I => \N__3234\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3237\,
            I => \N__3231\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3234\,
            I => \led_blink_inst.r_Count_2Z0Z_11\
        );

    \I__516\ : Odrv4
    port map (
            O => \N__3231\,
            I => \led_blink_inst.r_Count_2Z0Z_11\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__3226\,
            I => \N__3223\
        );

    \I__514\ : InMux
    port map (
            O => \N__3223\,
            I => \N__3220\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3220\,
            I => \N__3217\
        );

    \I__512\ : Odrv4
    port map (
            O => \N__3217\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_11\
        );

    \I__511\ : InMux
    port map (
            O => \N__3214\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_10\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__3211\,
            I => \N__3207\
        );

    \I__509\ : InMux
    port map (
            O => \N__3210\,
            I => \N__3204\
        );

    \I__508\ : InMux
    port map (
            O => \N__3207\,
            I => \N__3201\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3204\,
            I => \N__3198\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3201\,
            I => \led_blink_inst.r_Count_2Z0Z_12\
        );

    \I__505\ : Odrv4
    port map (
            O => \N__3198\,
            I => \led_blink_inst.r_Count_2Z0Z_12\
        );

    \I__504\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3190\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3190\,
            I => \N__3187\
        );

    \I__502\ : Span4Mux_v
    port map (
            O => \N__3187\,
            I => \N__3184\
        );

    \I__501\ : Odrv4
    port map (
            O => \N__3184\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_12\
        );

    \I__500\ : InMux
    port map (
            O => \N__3181\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_11\
        );

    \I__499\ : InMux
    port map (
            O => \N__3178\,
            I => \N__3175\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3175\,
            I => \led_blink_inst.o_LED_23_13\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__3172\,
            I => \led_blink_inst.o_LED_23_12_cascade_\
        );

    \I__496\ : InMux
    port map (
            O => \N__3169\,
            I => \N__3166\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3166\,
            I => \led_blink_inst.o_LED_23_15\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__3163\,
            I => \led_blink_inst.o_LED_23_21_cascade_\
        );

    \I__493\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3154\
        );

    \I__492\ : InMux
    port map (
            O => \N__3159\,
            I => \N__3154\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3154\,
            I => \N__3150\
        );

    \I__490\ : InMux
    port map (
            O => \N__3153\,
            I => \N__3147\
        );

    \I__489\ : Odrv4
    port map (
            O => \N__3150\,
            I => \led_blink_inst.r_Count_2Z0Z_1\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3147\,
            I => \led_blink_inst.r_Count_2Z0Z_1\
        );

    \I__487\ : CascadeMux
    port map (
            O => \N__3142\,
            I => \N__3138\
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__3141\,
            I => \N__3133\
        );

    \I__485\ : InMux
    port map (
            O => \N__3138\,
            I => \N__3126\
        );

    \I__484\ : InMux
    port map (
            O => \N__3137\,
            I => \N__3126\
        );

    \I__483\ : InMux
    port map (
            O => \N__3136\,
            I => \N__3126\
        );

    \I__482\ : InMux
    port map (
            O => \N__3133\,
            I => \N__3123\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3126\,
            I => \led_blink_inst.r_Count_2Z0Z_0\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3123\,
            I => \led_blink_inst.r_Count_2Z0Z_0\
        );

    \I__479\ : CascadeMux
    port map (
            O => \N__3118\,
            I => \N__3114\
        );

    \I__478\ : CascadeMux
    port map (
            O => \N__3117\,
            I => \N__3111\
        );

    \I__477\ : InMux
    port map (
            O => \N__3114\,
            I => \N__3108\
        );

    \I__476\ : InMux
    port map (
            O => \N__3111\,
            I => \N__3105\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__3108\,
            I => \led_blink_inst.r_Count_2Z0Z_2\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3105\,
            I => \led_blink_inst.r_Count_2Z0Z_2\
        );

    \I__473\ : InMux
    port map (
            O => \N__3100\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_1\
        );

    \I__472\ : InMux
    port map (
            O => \N__3097\,
            I => \N__3093\
        );

    \I__471\ : InMux
    port map (
            O => \N__3096\,
            I => \N__3090\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3093\,
            I => \led_blink_inst.r_Count_2Z0Z_3\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3090\,
            I => \led_blink_inst.r_Count_2Z0Z_3\
        );

    \I__468\ : InMux
    port map (
            O => \N__3085\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_2\
        );

    \I__467\ : InMux
    port map (
            O => \N__3082\,
            I => \N__3078\
        );

    \I__466\ : InMux
    port map (
            O => \N__3081\,
            I => \N__3075\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3078\,
            I => \led_blink_inst.r_Count_2Z0Z_4\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3075\,
            I => \led_blink_inst.r_Count_2Z0Z_4\
        );

    \I__463\ : InMux
    port map (
            O => \N__3070\,
            I => \N__3067\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3067\,
            I => \led_blink_inst.r_Count_2_RNO_0Z0Z_4\
        );

    \I__461\ : InMux
    port map (
            O => \N__3064\,
            I => \led_blink_inst.un2_r_Count_2_1_cry_3\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__3061\,
            I => \N__3058\
        );

    \I__459\ : InMux
    port map (
            O => \N__3058\,
            I => \N__3054\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__3057\,
            I => \N__3051\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3054\,
            I => \N__3048\
        );

    \I__456\ : InMux
    port map (
            O => \N__3051\,
            I => \N__3045\
        );

    \I__455\ : Odrv4
    port map (
            O => \N__3048\,
            I => \led_blink_inst.r_Count_1Z0Z_22\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3045\,
            I => \led_blink_inst.r_Count_1Z0Z_22\
        );

    \I__453\ : InMux
    port map (
            O => \N__3040\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_21\
        );

    \I__452\ : InMux
    port map (
            O => \N__3037\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_22\
        );

    \I__451\ : InMux
    port map (
            O => \N__3034\,
            I => \N__3031\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3031\,
            I => \N__3019\
        );

    \I__449\ : InMux
    port map (
            O => \N__3030\,
            I => \N__3010\
        );

    \I__448\ : InMux
    port map (
            O => \N__3029\,
            I => \N__3010\
        );

    \I__447\ : InMux
    port map (
            O => \N__3028\,
            I => \N__3010\
        );

    \I__446\ : InMux
    port map (
            O => \N__3027\,
            I => \N__3010\
        );

    \I__445\ : InMux
    port map (
            O => \N__3026\,
            I => \N__2999\
        );

    \I__444\ : InMux
    port map (
            O => \N__3025\,
            I => \N__2999\
        );

    \I__443\ : InMux
    port map (
            O => \N__3024\,
            I => \N__2999\
        );

    \I__442\ : InMux
    port map (
            O => \N__3023\,
            I => \N__2999\
        );

    \I__441\ : InMux
    port map (
            O => \N__3022\,
            I => \N__2999\
        );

    \I__440\ : Span4Mux_v
    port map (
            O => \N__3019\,
            I => \N__2992\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3010\,
            I => \N__2989\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2999\,
            I => \N__2986\
        );

    \I__437\ : InMux
    port map (
            O => \N__2998\,
            I => \N__2977\
        );

    \I__436\ : InMux
    port map (
            O => \N__2997\,
            I => \N__2977\
        );

    \I__435\ : InMux
    port map (
            O => \N__2996\,
            I => \N__2977\
        );

    \I__434\ : InMux
    port map (
            O => \N__2995\,
            I => \N__2977\
        );

    \I__433\ : Odrv4
    port map (
            O => \N__2992\,
            I => \led_blink_inst.o_LED_13_17\
        );

    \I__432\ : Odrv12
    port map (
            O => \N__2989\,
            I => \led_blink_inst.o_LED_13_17\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__2986\,
            I => \led_blink_inst.o_LED_13_17\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2977\,
            I => \led_blink_inst.o_LED_13_17\
        );

    \I__429\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2953\
        );

    \I__428\ : InMux
    port map (
            O => \N__2967\,
            I => \N__2944\
        );

    \I__427\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2944\
        );

    \I__426\ : InMux
    port map (
            O => \N__2965\,
            I => \N__2944\
        );

    \I__425\ : InMux
    port map (
            O => \N__2964\,
            I => \N__2944\
        );

    \I__424\ : InMux
    port map (
            O => \N__2963\,
            I => \N__2935\
        );

    \I__423\ : InMux
    port map (
            O => \N__2962\,
            I => \N__2935\
        );

    \I__422\ : InMux
    port map (
            O => \N__2961\,
            I => \N__2935\
        );

    \I__421\ : InMux
    port map (
            O => \N__2960\,
            I => \N__2935\
        );

    \I__420\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2926\
        );

    \I__419\ : InMux
    port map (
            O => \N__2958\,
            I => \N__2926\
        );

    \I__418\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2926\
        );

    \I__417\ : InMux
    port map (
            O => \N__2956\,
            I => \N__2926\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2953\,
            I => \led_blink_inst.o_LED_13_16\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2944\,
            I => \led_blink_inst.o_LED_13_16\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2935\,
            I => \led_blink_inst.o_LED_13_16\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2926\,
            I => \led_blink_inst.o_LED_13_16\
        );

    \I__412\ : CascadeMux
    port map (
            O => \N__2917\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_23_cascade_\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__2914\,
            I => \N__2903\
        );

    \I__410\ : CascadeMux
    port map (
            O => \N__2913\,
            I => \N__2900\
        );

    \I__409\ : CascadeMux
    port map (
            O => \N__2912\,
            I => \N__2897\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__2911\,
            I => \N__2892\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__2910\,
            I => \N__2887\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__2909\,
            I => \N__2884\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__2908\,
            I => \N__2881\
        );

    \I__404\ : InMux
    port map (
            O => \N__2907\,
            I => \N__2878\
        );

    \I__403\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2869\
        );

    \I__402\ : InMux
    port map (
            O => \N__2903\,
            I => \N__2869\
        );

    \I__401\ : InMux
    port map (
            O => \N__2900\,
            I => \N__2869\
        );

    \I__400\ : InMux
    port map (
            O => \N__2897\,
            I => \N__2869\
        );

    \I__399\ : InMux
    port map (
            O => \N__2896\,
            I => \N__2860\
        );

    \I__398\ : InMux
    port map (
            O => \N__2895\,
            I => \N__2860\
        );

    \I__397\ : InMux
    port map (
            O => \N__2892\,
            I => \N__2860\
        );

    \I__396\ : InMux
    port map (
            O => \N__2891\,
            I => \N__2860\
        );

    \I__395\ : InMux
    port map (
            O => \N__2890\,
            I => \N__2851\
        );

    \I__394\ : InMux
    port map (
            O => \N__2887\,
            I => \N__2851\
        );

    \I__393\ : InMux
    port map (
            O => \N__2884\,
            I => \N__2851\
        );

    \I__392\ : InMux
    port map (
            O => \N__2881\,
            I => \N__2851\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2878\,
            I => \led_blink_inst.o_LED_13_21\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__2869\,
            I => \led_blink_inst.o_LED_13_21\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2860\,
            I => \led_blink_inst.o_LED_13_21\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__2851\,
            I => \led_blink_inst.o_LED_13_21\
        );

    \I__387\ : CascadeMux
    port map (
            O => \N__2842\,
            I => \N__2839\
        );

    \I__386\ : InMux
    port map (
            O => \N__2839\,
            I => \N__2836\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2836\,
            I => \N__2832\
        );

    \I__384\ : InMux
    port map (
            O => \N__2835\,
            I => \N__2829\
        );

    \I__383\ : Odrv4
    port map (
            O => \N__2832\,
            I => \led_blink_inst.r_Count_1Z0Z_23\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2829\,
            I => \led_blink_inst.r_Count_1Z0Z_23\
        );

    \I__381\ : IoInMux
    port map (
            O => \N__2824\,
            I => \N__2821\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2821\,
            I => \N__2817\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__2820\,
            I => \N__2814\
        );

    \I__378\ : Span4Mux_s3_h
    port map (
            O => \N__2817\,
            I => \N__2811\
        );

    \I__377\ : InMux
    port map (
            O => \N__2814\,
            I => \N__2808\
        );

    \I__376\ : Odrv4
    port map (
            O => \N__2811\,
            I => \o_LED_2_c\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2808\,
            I => \o_LED_2_c\
        );

    \I__374\ : InMux
    port map (
            O => \N__2803\,
            I => \N__2800\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2800\,
            I => \N__2797\
        );

    \I__372\ : Odrv4
    port map (
            O => \N__2797\,
            I => \led_blink_inst.o_LED_23_14\
        );

    \I__371\ : CascadeMux
    port map (
            O => \N__2794\,
            I => \N__2790\
        );

    \I__370\ : CascadeMux
    port map (
            O => \N__2793\,
            I => \N__2787\
        );

    \I__369\ : InMux
    port map (
            O => \N__2790\,
            I => \N__2784\
        );

    \I__368\ : InMux
    port map (
            O => \N__2787\,
            I => \N__2781\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2784\,
            I => \led_blink_inst.r_Count_1Z0Z_14\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2781\,
            I => \led_blink_inst.r_Count_1Z0Z_14\
        );

    \I__365\ : InMux
    port map (
            O => \N__2776\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_13\
        );

    \I__364\ : CascadeMux
    port map (
            O => \N__2773\,
            I => \N__2769\
        );

    \I__363\ : InMux
    port map (
            O => \N__2772\,
            I => \N__2766\
        );

    \I__362\ : InMux
    port map (
            O => \N__2769\,
            I => \N__2763\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2766\,
            I => \led_blink_inst.r_Count_1Z0Z_15\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2763\,
            I => \led_blink_inst.r_Count_1Z0Z_15\
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__2758\,
            I => \N__2755\
        );

    \I__358\ : InMux
    port map (
            O => \N__2755\,
            I => \N__2752\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2752\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_15\
        );

    \I__356\ : InMux
    port map (
            O => \N__2749\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_14\
        );

    \I__355\ : InMux
    port map (
            O => \N__2746\,
            I => \N__2742\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__2745\,
            I => \N__2739\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2742\,
            I => \N__2736\
        );

    \I__352\ : InMux
    port map (
            O => \N__2739\,
            I => \N__2733\
        );

    \I__351\ : Odrv4
    port map (
            O => \N__2736\,
            I => \led_blink_inst.r_Count_1Z0Z_16\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2733\,
            I => \led_blink_inst.r_Count_1Z0Z_16\
        );

    \I__349\ : InMux
    port map (
            O => \N__2728\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_15\
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__2725\,
            I => \N__2721\
        );

    \I__347\ : InMux
    port map (
            O => \N__2724\,
            I => \N__2718\
        );

    \I__346\ : InMux
    port map (
            O => \N__2721\,
            I => \N__2715\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2718\,
            I => \led_blink_inst.r_Count_1Z0Z_17\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__2715\,
            I => \led_blink_inst.r_Count_1Z0Z_17\
        );

    \I__343\ : InMux
    port map (
            O => \N__2710\,
            I => \N__2707\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2707\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_17\
        );

    \I__341\ : InMux
    port map (
            O => \N__2704\,
            I => \bfn_8_9_0_\
        );

    \I__340\ : CascadeMux
    port map (
            O => \N__2701\,
            I => \N__2697\
        );

    \I__339\ : InMux
    port map (
            O => \N__2700\,
            I => \N__2694\
        );

    \I__338\ : InMux
    port map (
            O => \N__2697\,
            I => \N__2691\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2694\,
            I => \led_blink_inst.r_Count_1Z0Z_18\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2691\,
            I => \led_blink_inst.r_Count_1Z0Z_18\
        );

    \I__335\ : InMux
    port map (
            O => \N__2686\,
            I => \N__2683\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2683\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_18\
        );

    \I__333\ : InMux
    port map (
            O => \N__2680\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_17\
        );

    \I__332\ : CascadeMux
    port map (
            O => \N__2677\,
            I => \N__2673\
        );

    \I__331\ : InMux
    port map (
            O => \N__2676\,
            I => \N__2670\
        );

    \I__330\ : InMux
    port map (
            O => \N__2673\,
            I => \N__2667\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2670\,
            I => \led_blink_inst.r_Count_1Z0Z_19\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2667\,
            I => \led_blink_inst.r_Count_1Z0Z_19\
        );

    \I__327\ : InMux
    port map (
            O => \N__2662\,
            I => \N__2659\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2659\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_19\
        );

    \I__325\ : InMux
    port map (
            O => \N__2656\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_18\
        );

    \I__324\ : CascadeMux
    port map (
            O => \N__2653\,
            I => \N__2649\
        );

    \I__323\ : InMux
    port map (
            O => \N__2652\,
            I => \N__2646\
        );

    \I__322\ : InMux
    port map (
            O => \N__2649\,
            I => \N__2643\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2646\,
            I => \led_blink_inst.r_Count_1Z0Z_20\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2643\,
            I => \led_blink_inst.r_Count_1Z0Z_20\
        );

    \I__319\ : InMux
    port map (
            O => \N__2638\,
            I => \N__2635\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2635\,
            I => \N__2632\
        );

    \I__317\ : Span4Mux_h
    port map (
            O => \N__2632\,
            I => \N__2629\
        );

    \I__316\ : Odrv4
    port map (
            O => \N__2629\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_20\
        );

    \I__315\ : InMux
    port map (
            O => \N__2626\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_19\
        );

    \I__314\ : CascadeMux
    port map (
            O => \N__2623\,
            I => \N__2619\
        );

    \I__313\ : InMux
    port map (
            O => \N__2622\,
            I => \N__2616\
        );

    \I__312\ : InMux
    port map (
            O => \N__2619\,
            I => \N__2613\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2616\,
            I => \led_blink_inst.r_Count_1Z0Z_21\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2613\,
            I => \led_blink_inst.r_Count_1Z0Z_21\
        );

    \I__309\ : CascadeMux
    port map (
            O => \N__2608\,
            I => \N__2605\
        );

    \I__308\ : InMux
    port map (
            O => \N__2605\,
            I => \N__2602\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2602\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_21\
        );

    \I__306\ : InMux
    port map (
            O => \N__2599\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_20\
        );

    \I__305\ : InMux
    port map (
            O => \N__2596\,
            I => \N__2592\
        );

    \I__304\ : InMux
    port map (
            O => \N__2595\,
            I => \N__2589\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2592\,
            I => \led_blink_inst.r_Count_1Z0Z_6\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2589\,
            I => \led_blink_inst.r_Count_1Z0Z_6\
        );

    \I__301\ : InMux
    port map (
            O => \N__2584\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_5\
        );

    \I__300\ : InMux
    port map (
            O => \N__2581\,
            I => \N__2578\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2578\,
            I => \N__2575\
        );

    \I__298\ : Span4Mux_v
    port map (
            O => \N__2575\,
            I => \N__2571\
        );

    \I__297\ : InMux
    port map (
            O => \N__2574\,
            I => \N__2568\
        );

    \I__296\ : Odrv4
    port map (
            O => \N__2571\,
            I => \led_blink_inst.r_Count_1Z0Z_7\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2568\,
            I => \led_blink_inst.r_Count_1Z0Z_7\
        );

    \I__294\ : InMux
    port map (
            O => \N__2563\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_6\
        );

    \I__293\ : CascadeMux
    port map (
            O => \N__2560\,
            I => \N__2556\
        );

    \I__292\ : InMux
    port map (
            O => \N__2559\,
            I => \N__2553\
        );

    \I__291\ : InMux
    port map (
            O => \N__2556\,
            I => \N__2550\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2553\,
            I => \led_blink_inst.r_Count_1Z0Z_8\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2550\,
            I => \led_blink_inst.r_Count_1Z0Z_8\
        );

    \I__288\ : InMux
    port map (
            O => \N__2545\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_7\
        );

    \I__287\ : CascadeMux
    port map (
            O => \N__2542\,
            I => \N__2538\
        );

    \I__286\ : InMux
    port map (
            O => \N__2541\,
            I => \N__2535\
        );

    \I__285\ : InMux
    port map (
            O => \N__2538\,
            I => \N__2532\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2535\,
            I => \led_blink_inst.r_Count_1Z0Z_9\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2532\,
            I => \led_blink_inst.r_Count_1Z0Z_9\
        );

    \I__282\ : InMux
    port map (
            O => \N__2527\,
            I => \bfn_8_8_0_\
        );

    \I__281\ : InMux
    port map (
            O => \N__2524\,
            I => \N__2520\
        );

    \I__280\ : InMux
    port map (
            O => \N__2523\,
            I => \N__2517\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2520\,
            I => \led_blink_inst.r_Count_1Z0Z_10\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2517\,
            I => \led_blink_inst.r_Count_1Z0Z_10\
        );

    \I__277\ : CascadeMux
    port map (
            O => \N__2512\,
            I => \N__2509\
        );

    \I__276\ : InMux
    port map (
            O => \N__2509\,
            I => \N__2506\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2506\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_10\
        );

    \I__274\ : InMux
    port map (
            O => \N__2503\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_9\
        );

    \I__273\ : CascadeMux
    port map (
            O => \N__2500\,
            I => \N__2497\
        );

    \I__272\ : InMux
    port map (
            O => \N__2497\,
            I => \N__2493\
        );

    \I__271\ : InMux
    port map (
            O => \N__2496\,
            I => \N__2490\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2493\,
            I => \led_blink_inst.r_Count_1Z0Z_11\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2490\,
            I => \led_blink_inst.r_Count_1Z0Z_11\
        );

    \I__268\ : InMux
    port map (
            O => \N__2485\,
            I => \N__2482\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2482\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_11\
        );

    \I__266\ : InMux
    port map (
            O => \N__2479\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_10\
        );

    \I__265\ : CascadeMux
    port map (
            O => \N__2476\,
            I => \N__2472\
        );

    \I__264\ : InMux
    port map (
            O => \N__2475\,
            I => \N__2469\
        );

    \I__263\ : InMux
    port map (
            O => \N__2472\,
            I => \N__2466\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2469\,
            I => \led_blink_inst.r_Count_1Z0Z_12\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2466\,
            I => \led_blink_inst.r_Count_1Z0Z_12\
        );

    \I__260\ : InMux
    port map (
            O => \N__2461\,
            I => \N__2458\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__2458\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_12\
        );

    \I__258\ : InMux
    port map (
            O => \N__2455\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_11\
        );

    \I__257\ : CascadeMux
    port map (
            O => \N__2452\,
            I => \N__2448\
        );

    \I__256\ : InMux
    port map (
            O => \N__2451\,
            I => \N__2445\
        );

    \I__255\ : InMux
    port map (
            O => \N__2448\,
            I => \N__2442\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2445\,
            I => \led_blink_inst.r_Count_1Z0Z_13\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2442\,
            I => \led_blink_inst.r_Count_1Z0Z_13\
        );

    \I__252\ : CascadeMux
    port map (
            O => \N__2437\,
            I => \N__2434\
        );

    \I__251\ : InMux
    port map (
            O => \N__2434\,
            I => \N__2431\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2431\,
            I => \N__2428\
        );

    \I__249\ : Odrv4
    port map (
            O => \N__2428\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_13\
        );

    \I__248\ : InMux
    port map (
            O => \N__2425\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_12\
        );

    \I__247\ : InMux
    port map (
            O => \N__2422\,
            I => \N__2417\
        );

    \I__246\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2414\
        );

    \I__245\ : InMux
    port map (
            O => \N__2420\,
            I => \N__2411\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__2417\,
            I => \led_blink_inst.r_Count_1Z0Z_1\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2414\,
            I => \led_blink_inst.r_Count_1Z0Z_1\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__2411\,
            I => \led_blink_inst.r_Count_1Z0Z_1\
        );

    \I__241\ : CascadeMux
    port map (
            O => \N__2404\,
            I => \N__2398\
        );

    \I__240\ : InMux
    port map (
            O => \N__2403\,
            I => \N__2395\
        );

    \I__239\ : InMux
    port map (
            O => \N__2402\,
            I => \N__2392\
        );

    \I__238\ : InMux
    port map (
            O => \N__2401\,
            I => \N__2389\
        );

    \I__237\ : InMux
    port map (
            O => \N__2398\,
            I => \N__2386\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2395\,
            I => \led_blink_inst.r_Count_1Z0Z_0\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__2392\,
            I => \led_blink_inst.r_Count_1Z0Z_0\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2389\,
            I => \led_blink_inst.r_Count_1Z0Z_0\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2386\,
            I => \led_blink_inst.r_Count_1Z0Z_0\
        );

    \I__232\ : CascadeMux
    port map (
            O => \N__2377\,
            I => \N__2374\
        );

    \I__231\ : InMux
    port map (
            O => \N__2374\,
            I => \N__2370\
        );

    \I__230\ : InMux
    port map (
            O => \N__2373\,
            I => \N__2367\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2370\,
            I => \led_blink_inst.r_Count_1Z0Z_2\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__2367\,
            I => \led_blink_inst.r_Count_1Z0Z_2\
        );

    \I__227\ : InMux
    port map (
            O => \N__2362\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_1\
        );

    \I__226\ : InMux
    port map (
            O => \N__2359\,
            I => \N__2355\
        );

    \I__225\ : InMux
    port map (
            O => \N__2358\,
            I => \N__2352\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2355\,
            I => \led_blink_inst.r_Count_1Z0Z_3\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__2352\,
            I => \led_blink_inst.r_Count_1Z0Z_3\
        );

    \I__222\ : InMux
    port map (
            O => \N__2347\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_2\
        );

    \I__221\ : CascadeMux
    port map (
            O => \N__2344\,
            I => \N__2340\
        );

    \I__220\ : InMux
    port map (
            O => \N__2343\,
            I => \N__2337\
        );

    \I__219\ : InMux
    port map (
            O => \N__2340\,
            I => \N__2334\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__2337\,
            I => \led_blink_inst.r_Count_1Z0Z_4\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__2334\,
            I => \led_blink_inst.r_Count_1Z0Z_4\
        );

    \I__216\ : InMux
    port map (
            O => \N__2329\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_3\
        );

    \I__215\ : InMux
    port map (
            O => \N__2326\,
            I => \N__2322\
        );

    \I__214\ : InMux
    port map (
            O => \N__2325\,
            I => \N__2319\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__2322\,
            I => \led_blink_inst.r_Count_1Z0Z_5\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__2319\,
            I => \led_blink_inst.r_Count_1Z0Z_5\
        );

    \I__211\ : InMux
    port map (
            O => \N__2314\,
            I => \N__2311\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__2311\,
            I => \led_blink_inst.r_Count_1_RNO_0Z0Z_5\
        );

    \I__209\ : InMux
    port map (
            O => \N__2308\,
            I => \led_blink_inst.un3_r_Count_1_1_cry_4\
        );

    \I__208\ : CascadeMux
    port map (
            O => \N__2305\,
            I => \led_blink_inst.o_LED_23_16_cascade_\
        );

    \I__207\ : InMux
    port map (
            O => \N__2302\,
            I => \N__2299\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__2299\,
            I => \led_blink_inst.o_LED_13_15\
        );

    \I__205\ : InMux
    port map (
            O => \N__2296\,
            I => \N__2293\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__2293\,
            I => \led_blink_inst.o_LED_13_13\
        );

    \I__203\ : CascadeMux
    port map (
            O => \N__2290\,
            I => \led_blink_inst.o_LED_13_14_cascade_\
        );

    \I__202\ : InMux
    port map (
            O => \N__2287\,
            I => \N__2284\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__2284\,
            I => \led_blink_inst.o_LED_13_12\
        );

    \I__200\ : CascadeMux
    port map (
            O => \N__2281\,
            I => \led_blink_inst.o_LED_13_21_cascade_\
        );

    \I__199\ : CascadeMux
    port map (
            O => \N__2278\,
            I => \led_blink_inst.o_LED_13_16_cascade_\
        );

    \I__198\ : IoInMux
    port map (
            O => \N__2275\,
            I => \N__2272\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__2272\,
            I => \N__2269\
        );

    \I__196\ : IoSpan4Mux
    port map (
            O => \N__2269\,
            I => \N__2266\
        );

    \I__195\ : Span4Mux_s3_h
    port map (
            O => \N__2266\,
            I => \N__2262\
        );

    \I__194\ : InMux
    port map (
            O => \N__2265\,
            I => \N__2259\
        );

    \I__193\ : Odrv4
    port map (
            O => \N__2262\,
            I => \o_LED_1_c\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__2259\,
            I => \o_LED_1_c\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \led_blink_inst.un3_r_Count_1_1_cry_8\,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \led_blink_inst.un3_r_Count_1_1_cry_16\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \led_blink_inst.un2_r_Count_4_1_cry_8\,
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \led_blink_inst.un2_r_Count_4_1_cry_16\,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_12_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_3_0_\
        );

    \IN_MUX_bfv_12_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \led_blink_inst.un2_r_Count_3_1_cry_8\,
            carryinitout => \bfn_12_4_0_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \led_blink_inst.un2_r_Count_3_1_cry_16\,
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \led_blink_inst.un2_r_Count_2_1_cry_8\,
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \led_blink_inst.un2_r_Count_2_1_cry_16\,
            carryinitout => \bfn_9_8_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNIVTTA_13_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2772\,
            in1 => \N__2451\,
            in2 => \N__2701\,
            in3 => \N__2724\,
            lcout => \led_blink_inst.o_LED_13_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNIJ5RV_16_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2746\,
            in1 => \N__2343\,
            in2 => \N__3061\,
            in3 => \N__2401\,
            lcout => \led_blink_inst.o_LED_13_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__2996\,
            in1 => \N__2957\,
            in2 => \N__2909\,
            in3 => \N__2402\,
            lcout => \led_blink_inst.r_Count_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNILPMK1_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2421\,
            in1 => \N__2596\,
            in2 => \N__2377\,
            in3 => \N__2559\,
            lcout => \led_blink_inst.o_LED_13_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNICN8A1_14_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2581\,
            in1 => \N__2359\,
            in2 => \N__2794\,
            in3 => \N__2541\,
            lcout => \led_blink_inst.o_LED_13_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.o_LED_1_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__2995\,
            in1 => \N__2265\,
            in2 => \N__2908\,
            in3 => \N__2956\,
            lcout => \o_LED_1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_5_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2998\,
            in1 => \N__2959\,
            in2 => \N__2910\,
            in3 => \N__2314\,
            lcout => \led_blink_inst.r_Count_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_15_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__2958\,
            in1 => \N__2997\,
            in2 => \N__2758\,
            in3 => \N__2890\,
            lcout => \led_blink_inst.r_Count_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNIVMBL_10_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2524\,
            in1 => \N__2326\,
            in2 => \N__2500\,
            in3 => \N__2475\,
            lcout => OPEN,
            ltout => \led_blink_inst.o_LED_13_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNIV59V3_10_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2302\,
            in1 => \N__2296\,
            in2 => \N__2290\,
            in3 => \N__2287\,
            lcout => \led_blink_inst.o_LED_13_21\,
            ltout => \led_blink_inst.o_LED_13_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_20_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2963\,
            in1 => \N__3026\,
            in2 => \N__2281\,
            in3 => \N__2638\,
            lcout => \led_blink_inst.r_Count_1Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNIOP0B_23_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2622\,
            in1 => \N__2652\,
            in2 => \N__2842\,
            in3 => \N__2676\,
            lcout => \led_blink_inst.o_LED_13_16\,
            ltout => \led_blink_inst.o_LED_13_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_11_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2891\,
            in1 => \N__3023\,
            in2 => \N__2278\,
            in3 => \N__2485\,
            lcout => \led_blink_inst.r_Count_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_13_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3025\,
            in1 => \N__2962\,
            in2 => \N__2437\,
            in3 => \N__2896\,
            lcout => \led_blink_inst.r_Count_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_12_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2961\,
            in1 => \N__3024\,
            in2 => \N__2911\,
            in3 => \N__2461\,
            lcout => \led_blink_inst.r_Count_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_10_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3022\,
            in1 => \N__2960\,
            in2 => \N__2512\,
            in3 => \N__2895\,
            lcout => \led_blink_inst.r_Count_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_18_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3028\,
            in1 => \N__2965\,
            in2 => \N__2913\,
            in3 => \N__2686\,
            lcout => \led_blink_inst.r_Count_1Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_17_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3027\,
            in1 => \N__2964\,
            in2 => \N__2912\,
            in3 => \N__2710\,
            lcout => \led_blink_inst.r_Count_1Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_19_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3029\,
            in1 => \N__2966\,
            in2 => \N__2914\,
            in3 => \N__2662\,
            lcout => \led_blink_inst.r_Count_1Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_21_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__2967\,
            in1 => \N__3030\,
            in2 => \N__2608\,
            in3 => \N__2906\,
            lcout => \led_blink_inst.r_Count_1Z0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNI1EOR_18_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3393\,
            in1 => \N__3426\,
            in2 => \N__3604\,
            in3 => \N__3453\,
            lcout => \led_blink_inst.o_LED_23_16\,
            ltout => \led_blink_inst.o_LED_23_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_12_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__3193\,
            in1 => \N__3791\,
            in2 => \N__2305\,
            in3 => \N__3655\,
            lcout => \led_blink_inst.r_Count_2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNIOJCA1_10_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3301\,
            in1 => \N__3082\,
            in2 => \N__3244\,
            in3 => \N__3270\,
            lcout => \led_blink_inst.o_LED_23_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNIV9MR_12_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3562\,
            in1 => \N__3519\,
            in2 => \N__3211\,
            in3 => \N__3489\,
            lcout => \led_blink_inst.o_LED_23_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_17_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3794\,
            in1 => \N__3729\,
            in2 => \N__3475\,
            in3 => \N__3660\,
            lcout => \led_blink_inst.r_Count_2Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2403\,
            in2 => \_gnd_net_\,
            in3 => \N__2422\,
            lcout => \led_blink_inst.r_Count_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_20_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3797\,
            in1 => \N__3732\,
            in2 => \N__3379\,
            in3 => \N__3665\,
            lcout => \led_blink_inst.r_Count_2Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_19_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3796\,
            in1 => \N__3731\,
            in2 => \N__3412\,
            in3 => \N__3664\,
            lcout => \led_blink_inst.r_Count_2Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_18_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3730\,
            in1 => \N__3795\,
            in2 => \N__3672\,
            in3 => \N__3439\,
            lcout => \led_blink_inst.r_Count_2Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_10_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3792\,
            in1 => \N__3727\,
            in2 => \N__3256\,
            in3 => \N__3656\,
            lcout => \led_blink_inst.r_Count_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_14_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3728\,
            in1 => \N__3793\,
            in2 => \N__3671\,
            in3 => \N__3550\,
            lcout => \led_blink_inst.r_Count_2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.un3_r_Count_1_1_cry_1_c_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2420\,
            in2 => \N__2404\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_2_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2373\,
            in2 => \_gnd_net_\,
            in3 => \N__2362\,
            lcout => \led_blink_inst.r_Count_1Z0Z_2\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_1\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_2\,
            clk => \N__4932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_3_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2358\,
            in2 => \_gnd_net_\,
            in3 => \N__2347\,
            lcout => \led_blink_inst.r_Count_1Z0Z_3\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_2\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_3\,
            clk => \N__4932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_4_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2344\,
            in3 => \N__2329\,
            lcout => \led_blink_inst.r_Count_1Z0Z_4\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_3\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_4\,
            clk => \N__4932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_5_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2325\,
            in2 => \_gnd_net_\,
            in3 => \N__2308\,
            lcout => \led_blink_inst.r_Count_1_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_4\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_6_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2595\,
            in2 => \_gnd_net_\,
            in3 => \N__2584\,
            lcout => \led_blink_inst.r_Count_1Z0Z_6\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_5\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_6\,
            clk => \N__4932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_7_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2574\,
            in2 => \_gnd_net_\,
            in3 => \N__2563\,
            lcout => \led_blink_inst.r_Count_1Z0Z_7\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_6\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_7\,
            clk => \N__4932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_8_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2560\,
            in3 => \N__2545\,
            lcout => \led_blink_inst.r_Count_1Z0Z_8\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_7\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_8\,
            clk => \N__4932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_9_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2542\,
            in3 => \N__2527\,
            lcout => \led_blink_inst.r_Count_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_9\,
            clk => \N__4928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_10_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2523\,
            in2 => \_gnd_net_\,
            in3 => \N__2503\,
            lcout => \led_blink_inst.r_Count_1_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_9\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_11_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2496\,
            in2 => \_gnd_net_\,
            in3 => \N__2479\,
            lcout => \led_blink_inst.r_Count_1_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_10\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_12_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2476\,
            in3 => \N__2455\,
            lcout => \led_blink_inst.r_Count_1_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_11\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_13_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2452\,
            in3 => \N__2425\,
            lcout => \led_blink_inst.r_Count_1_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_12\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_14_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2793\,
            in3 => \N__2776\,
            lcout => \led_blink_inst.r_Count_1Z0Z_14\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_13\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_14\,
            clk => \N__4928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_15_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2773\,
            in3 => \N__2749\,
            lcout => \led_blink_inst.r_Count_1_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_14\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_16_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2745\,
            in3 => \N__2728\,
            lcout => \led_blink_inst.r_Count_1Z0Z_16\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_15\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_16\,
            clk => \N__4928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_17_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2725\,
            in3 => \N__2704\,
            lcout => \led_blink_inst.r_Count_1_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_18_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2700\,
            in2 => \_gnd_net_\,
            in3 => \N__2680\,
            lcout => \led_blink_inst.r_Count_1_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_17\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_19_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2677\,
            in3 => \N__2656\,
            lcout => \led_blink_inst.r_Count_1_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_18\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_20_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2653\,
            in3 => \N__2626\,
            lcout => \led_blink_inst.r_Count_1_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_19\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_21_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2623\,
            in3 => \N__2599\,
            lcout => \led_blink_inst.r_Count_1_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_20\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_22_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3057\,
            in3 => \N__3040\,
            lcout => \led_blink_inst.r_Count_1Z0Z_22\,
            ltout => OPEN,
            carryin => \led_blink_inst.un3_r_Count_1_1_cry_21\,
            carryout => \led_blink_inst.un3_r_Count_1_1_cry_22\,
            clk => \N__4933\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_RNO_0_23_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2835\,
            in2 => \_gnd_net_\,
            in3 => \N__3037\,
            lcout => OPEN,
            ltout => \led_blink_inst.r_Count_1_RNO_0Z0Z_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_1_23_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3034\,
            in1 => \N__2968\,
            in2 => \N__2917\,
            in3 => \N__2907\,
            lcout => \led_blink_inst.r_Count_1Z0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4933\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_11_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3725\,
            in1 => \N__3789\,
            in2 => \N__3226\,
            in3 => \N__3651\,
            lcout => \led_blink_inst.r_Count_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_16_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3790\,
            in1 => \N__3726\,
            in2 => \N__3670\,
            in3 => \N__3505\,
            lcout => \led_blink_inst.r_Count_2Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.o_LED_2_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__3724\,
            in1 => \N__3788\,
            in2 => \N__2820\,
            in3 => \N__3650\,
            lcout => \o_LED_2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_1_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3160\,
            in1 => \_gnd_net_\,
            in2 => \N__3142\,
            in3 => \_gnd_net_\,
            lcout => \led_blink_inst.r_Count_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNI0SCA1_13_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3349\,
            in1 => \N__3316\,
            in2 => \N__3583\,
            in3 => \N__3541\,
            lcout => \led_blink_inst.o_LED_23_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNI7SOH1_23_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3364\,
            in1 => \N__3097\,
            in2 => \N__3118\,
            in3 => \N__3817\,
            lcout => OPEN,
            ltout => \led_blink_inst.o_LED_23_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNIUL825_10_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2803\,
            in1 => \N__3178\,
            in2 => \N__3172\,
            in3 => \N__3169\,
            lcout => \led_blink_inst.o_LED_23_21\,
            ltout => \led_blink_inst.o_LED_23_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_9_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3787\,
            in1 => \N__3723\,
            in2 => \N__3163\,
            in3 => \N__3283\,
            lcout => \led_blink_inst.r_Count_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_4_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3722\,
            in1 => \N__3786\,
            in2 => \N__3669\,
            in3 => \N__3070\,
            lcout => \led_blink_inst.r_Count_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_0_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__3137\,
            in1 => \N__3721\,
            in2 => \N__3801\,
            in3 => \N__3646\,
            lcout => \led_blink_inst.r_Count_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNI3OOH1_21_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3333\,
            in1 => \N__3136\,
            in2 => \N__3847\,
            in3 => \N__3159\,
            lcout => \led_blink_inst.o_LED_23_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.un2_r_Count_2_1_cry_1_c_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3153\,
            in2 => \N__3141\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_2_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3117\,
            in3 => \N__3100\,
            lcout => \led_blink_inst.r_Count_2Z0Z_2\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_1\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_2\,
            clk => \N__4938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_3_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3096\,
            in2 => \_gnd_net_\,
            in3 => \N__3085\,
            lcout => \led_blink_inst.r_Count_2Z0Z_3\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_2\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_3\,
            clk => \N__4938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_4_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3081\,
            in2 => \_gnd_net_\,
            in3 => \N__3064\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_3\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_5_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3363\,
            in2 => \_gnd_net_\,
            in3 => \N__3352\,
            lcout => \led_blink_inst.r_Count_2Z0Z_5\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_4\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_5\,
            clk => \N__4938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_6_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3348\,
            in2 => \_gnd_net_\,
            in3 => \N__3337\,
            lcout => \led_blink_inst.r_Count_2Z0Z_6\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_5\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_6\,
            clk => \N__4938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_7_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3334\,
            in3 => \N__3319\,
            lcout => \led_blink_inst.r_Count_2Z0Z_7\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_6\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_7\,
            clk => \N__4938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_8_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3315\,
            in2 => \_gnd_net_\,
            in3 => \N__3304\,
            lcout => \led_blink_inst.r_Count_2Z0Z_8\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_7\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_8\,
            clk => \N__4938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_9_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3300\,
            in2 => \_gnd_net_\,
            in3 => \N__3274\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_10_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3271\,
            in3 => \N__3247\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_9\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_11_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3243\,
            in2 => \_gnd_net_\,
            in3 => \N__3214\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_10\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_12_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3210\,
            in2 => \_gnd_net_\,
            in3 => \N__3181\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_11\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_13_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3576\,
            in2 => \_gnd_net_\,
            in3 => \N__3565\,
            lcout => \led_blink_inst.r_Count_2Z0Z_13\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_12\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_13\,
            clk => \N__4935\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_14_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3561\,
            in2 => \_gnd_net_\,
            in3 => \N__3544\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_13\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_15_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3540\,
            in3 => \N__3523\,
            lcout => \led_blink_inst.r_Count_2Z0Z_15\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_14\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_15\,
            clk => \N__4935\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_16_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3520\,
            in2 => \_gnd_net_\,
            in3 => \N__3496\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_15\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_17_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3493\,
            in3 => \N__3460\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_18_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3457\,
            in3 => \N__3430\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_17\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_19_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3427\,
            in2 => \_gnd_net_\,
            in3 => \N__3400\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_18\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_20_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3397\,
            in3 => \N__3367\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_19\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_21_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3843\,
            in3 => \N__3826\,
            lcout => \led_blink_inst.r_Count_2Z0Z_21\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_20\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_21\,
            clk => \N__4931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_RNO_0_22_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3594\,
            in2 => \_gnd_net_\,
            in3 => \N__3823\,
            lcout => \led_blink_inst.r_Count_2_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_2_1_cry_21\,
            carryout => \led_blink_inst.un2_r_Count_2_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_23_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3816\,
            in2 => \_gnd_net_\,
            in3 => \N__3820\,
            lcout => \led_blink_inst.r_Count_2Z0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_2_22_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3802\,
            in1 => \N__3739\,
            in2 => \N__3682\,
            in3 => \N__3673\,
            lcout => \led_blink_inst.r_Count_2Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNI527P1_11_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4297\,
            in1 => \N__4113\,
            in2 => \N__4435\,
            in3 => \N__4266\,
            lcout => \led_blink_inst.o_LED_33_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_8_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4038\,
            in1 => \N__3994\,
            in2 => \N__4171\,
            in3 => \N__3954\,
            lcout => \led_blink_inst.r_Count_3Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_7_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4037\,
            in1 => \N__3993\,
            in2 => \N__3958\,
            in3 => \N__4195\,
            lcout => \led_blink_inst.r_Count_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNIHE7P1_10_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4210\,
            in1 => \N__4249\,
            in2 => \N__4462\,
            in3 => \N__4185\,
            lcout => \led_blink_inst.o_LED_33_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_5_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4036\,
            in1 => \N__3992\,
            in2 => \N__3957\,
            in3 => \N__4237\,
            lcout => \led_blink_inst.r_Count_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_1_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__4098\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4114\,
            lcout => \led_blink_inst.r_Count_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNIU40L1_23_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4338\,
            in1 => \N__4228\,
            in2 => \N__4507\,
            in3 => \N__4096\,
            lcout => \led_blink_inst.o_LED_33_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNIK2NG1_14_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4375\,
            in1 => \N__4282\,
            in2 => \N__4591\,
            in3 => \N__4356\,
            lcout => OPEN,
            ltout => \led_blink_inst.o_LED_33_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNIEFLF6_10_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3892\,
            in1 => \N__3883\,
            in2 => \N__3877\,
            in3 => \N__4048\,
            lcout => \led_blink_inst.o_LED_33_21\,
            ltout => \led_blink_inst.o_LED_33_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.o_LED_3_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__3867\,
            in1 => \N__4023\,
            in2 => \N__3874\,
            in3 => \N__3986\,
            lcout => \o_LED_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4947\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_10_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3988\,
            in1 => \N__4027\,
            in2 => \N__3955\,
            in3 => \N__4444\,
            lcout => \led_blink_inst.r_Count_3Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4947\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNIEUOG1_12_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4569\,
            in1 => \N__4413\,
            in2 => \N__4528\,
            in3 => \N__4155\,
            lcout => \led_blink_inst.o_LED_33_16\,
            ltout => \led_blink_inst.o_LED_33_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_13_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3941\,
            in1 => \N__4028\,
            in2 => \N__3850\,
            in3 => \N__4384\,
            lcout => \led_blink_inst.r_Count_3Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4947\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_0_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__4097\,
            in1 => \N__3987\,
            in2 => \N__4039\,
            in3 => \N__3942\,
            lcout => \led_blink_inst.r_Count_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4947\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_21_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3991\,
            in1 => \N__4042\,
            in2 => \N__3956\,
            in3 => \N__4537\,
            lcout => \led_blink_inst.r_Count_3Z0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_17_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4040\,
            in1 => \N__3989\,
            in2 => \N__4309\,
            in3 => \N__3946\,
            lcout => \led_blink_inst.r_Count_3Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNI4SFC1_13_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4320\,
            in1 => \N__4396\,
            in2 => \N__4552\,
            in3 => \N__4617\,
            lcout => \led_blink_inst.o_LED_33_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_18_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4041\,
            in1 => \N__3990\,
            in2 => \N__4603\,
            in3 => \N__3947\,
            lcout => \led_blink_inst.r_Count_3Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.un2_r_Count_4_1_cry_1_c_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5170\,
            in2 => \N__5136\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_2_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5244\,
            in2 => \_gnd_net_\,
            in3 => \N__3907\,
            lcout => \led_blink_inst.r_Count_4Z0Z_2\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_1\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_2\,
            clk => \N__4942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_3_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4629\,
            in2 => \_gnd_net_\,
            in3 => \N__3904\,
            lcout => \led_blink_inst.r_Count_4Z0Z_3\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_2\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_3\,
            clk => \N__4942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNO_0_4_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4761\,
            in2 => \_gnd_net_\,
            in3 => \N__3901\,
            lcout => \led_blink_inst.r_Count_4_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_3\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_5_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4705\,
            in3 => \N__3898\,
            lcout => \led_blink_inst.r_Count_4Z0Z_5\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_4\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_5\,
            clk => \N__4942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNO_0_6_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4800\,
            in2 => \_gnd_net_\,
            in3 => \N__3895\,
            lcout => \led_blink_inst.r_Count_4_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_5\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNO_0_7_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4773\,
            in2 => \_gnd_net_\,
            in3 => \N__4075\,
            lcout => \led_blink_inst.r_Count_4_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_6\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_8_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4750\,
            in3 => \N__4072\,
            lcout => \led_blink_inst.r_Count_4Z0Z_8\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_7\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_8\,
            clk => \N__4942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNO_0_9_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4788\,
            in2 => \_gnd_net_\,
            in3 => \N__4069\,
            lcout => \led_blink_inst.r_Count_4_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_10_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4734\,
            in2 => \_gnd_net_\,
            in3 => \N__4066\,
            lcout => \led_blink_inst.r_Count_4Z0Z_10\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_9\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_10\,
            clk => \N__4940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_11_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5256\,
            in2 => \_gnd_net_\,
            in3 => \N__4063\,
            lcout => \led_blink_inst.r_Count_4Z0Z_11\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_10\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_11\,
            clk => \N__4940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNO_0_12_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4870\,
            in2 => \_gnd_net_\,
            in3 => \N__4060\,
            lcout => \led_blink_inst.r_Count_4_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_11\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_13_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4722\,
            in3 => \N__4057\,
            lcout => \led_blink_inst.r_Count_4Z0Z_13\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_12\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_13\,
            clk => \N__4940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_14_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4668\,
            in2 => \_gnd_net_\,
            in3 => \N__4054\,
            lcout => \led_blink_inst.r_Count_4Z0Z_14\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_13\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_14\,
            clk => \N__4940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_15_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5215\,
            in3 => \N__4051\,
            lcout => \led_blink_inst.r_Count_4Z0Z_15\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_14\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_15\,
            clk => \N__4940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNO_0_16_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4855\,
            in3 => \N__4138\,
            lcout => \led_blink_inst.r_Count_4_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_15\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNO_0_17_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4839\,
            in2 => \_gnd_net_\,
            in3 => \N__4135\,
            lcout => \led_blink_inst.r_Count_4_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_18_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5232\,
            in3 => \N__4132\,
            lcout => \led_blink_inst.r_Count_4Z0Z_18\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_17\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_18\,
            clk => \N__4936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_19_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5191\,
            in3 => \N__4129\,
            lcout => \led_blink_inst.r_Count_4Z0Z_19\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_18\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_19\,
            clk => \N__4936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNO_0_20_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4825\,
            in2 => \_gnd_net_\,
            in3 => \N__4126\,
            lcout => \led_blink_inst.r_Count_4_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_19\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_21_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4644\,
            in2 => \_gnd_net_\,
            in3 => \N__4123\,
            lcout => \led_blink_inst.r_Count_4Z0Z_21\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_20\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_21\,
            clk => \N__4936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_22_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5151\,
            in2 => \_gnd_net_\,
            in3 => \N__4120\,
            lcout => \led_blink_inst.r_Count_4Z0Z_22\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_4_1_cry_21\,
            carryout => \led_blink_inst.un2_r_Count_4_1_cry_22\,
            clk => \N__4936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_23_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4657\,
            in2 => \_gnd_net_\,
            in3 => \N__4117\,
            lcout => \led_blink_inst.r_Count_4Z0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.un2_r_Count_3_1_cry_1_c_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4112\,
            in2 => \N__4099\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_3_0_\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_2_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4296\,
            in2 => \_gnd_net_\,
            in3 => \N__4285\,
            lcout => \led_blink_inst.r_Count_3Z0Z_2\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_1\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_2\,
            clk => \N__4951\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_3_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4281\,
            in2 => \_gnd_net_\,
            in3 => \N__4270\,
            lcout => \led_blink_inst.r_Count_3Z0Z_3\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_2\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_3\,
            clk => \N__4951\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_4_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4267\,
            in3 => \N__4252\,
            lcout => \led_blink_inst.r_Count_3Z0Z_4\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_3\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_4\,
            clk => \N__4951\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNO_0_5_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4248\,
            in2 => \_gnd_net_\,
            in3 => \N__4231\,
            lcout => \led_blink_inst.r_Count_3_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_4\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_6_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4224\,
            in2 => \_gnd_net_\,
            in3 => \N__4213\,
            lcout => \led_blink_inst.r_Count_3Z0Z_6\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_5\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_6\,
            clk => \N__4951\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNO_0_7_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4206\,
            in2 => \_gnd_net_\,
            in3 => \N__4189\,
            lcout => \led_blink_inst.r_Count_3_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_6\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNO_0_8_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4186\,
            in3 => \N__4159\,
            lcout => \led_blink_inst.r_Count_3_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_7\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_9_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4156\,
            in3 => \N__4141\,
            lcout => \led_blink_inst.r_Count_3Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_4_0_\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_9\,
            clk => \N__4950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNO_0_10_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4461\,
            in3 => \N__4438\,
            lcout => \led_blink_inst.r_Count_3_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_9\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_11_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4434\,
            in3 => \N__4417\,
            lcout => \led_blink_inst.r_Count_3Z0Z_11\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_10\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_11\,
            clk => \N__4950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_12_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4414\,
            in3 => \N__4399\,
            lcout => \led_blink_inst.r_Count_3Z0Z_12\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_11\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_12\,
            clk => \N__4950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNO_0_13_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4395\,
            in2 => \_gnd_net_\,
            in3 => \N__4378\,
            lcout => \led_blink_inst.r_Count_3_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_12\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_14_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4371\,
            in2 => \_gnd_net_\,
            in3 => \N__4360\,
            lcout => \led_blink_inst.r_Count_3Z0Z_14\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_13\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_14\,
            clk => \N__4950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_15_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4357\,
            in3 => \N__4342\,
            lcout => \led_blink_inst.r_Count_3Z0Z_15\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_14\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_15\,
            clk => \N__4950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_16_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4339\,
            in3 => \N__4324\,
            lcout => \led_blink_inst.r_Count_3Z0Z_16\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_15\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_16\,
            clk => \N__4950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNO_0_17_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4321\,
            in2 => \_gnd_net_\,
            in3 => \N__4300\,
            lcout => \led_blink_inst.r_Count_3_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNO_0_18_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4618\,
            in3 => \N__4594\,
            lcout => \led_blink_inst.r_Count_3_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_17\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_19_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4590\,
            in3 => \N__4573\,
            lcout => \led_blink_inst.r_Count_3Z0Z_19\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_18\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_19\,
            clk => \N__4948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_20_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4570\,
            in3 => \N__4555\,
            lcout => \led_blink_inst.r_Count_3Z0Z_20\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_19\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_20\,
            clk => \N__4948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_RNO_0_21_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4551\,
            in2 => \_gnd_net_\,
            in3 => \N__4531\,
            lcout => \led_blink_inst.r_Count_3_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_20\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_22_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4527\,
            in2 => \_gnd_net_\,
            in3 => \N__4513\,
            lcout => \led_blink_inst.r_Count_3Z0Z_22\,
            ltout => OPEN,
            carryin => \led_blink_inst.un2_r_Count_3_1_cry_21\,
            carryout => \led_blink_inst.un2_r_Count_3_1_cry_22\,
            clk => \N__4948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_3_23_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4503\,
            in2 => \_gnd_net_\,
            in3 => \N__4510\,
            lcout => \led_blink_inst.r_Count_3Z0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_4_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4992\,
            in1 => \N__5037\,
            in2 => \N__4489\,
            in3 => \N__5087\,
            lcout => \led_blink_inst.r_Count_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_7_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5039\,
            in1 => \N__4989\,
            in2 => \N__5091\,
            in3 => \N__4477\,
            lcout => \led_blink_inst.r_Count_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_6_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4993\,
            in1 => \N__5038\,
            in2 => \N__4471\,
            in3 => \N__5088\,
            lcout => \led_blink_inst.r_Count_4Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_9_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5040\,
            in1 => \N__4990\,
            in2 => \N__5092\,
            in3 => \N__4807\,
            lcout => \led_blink_inst.r_Count_4Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNIA7S1_4_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4801\,
            in1 => \N__4789\,
            in2 => \N__4777\,
            in3 => \N__4762\,
            lcout => \led_blink_inst.o_LED_43_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNI2IHV_5_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4749\,
            in1 => \N__4735\,
            in2 => \N__4723\,
            in3 => \N__4704\,
            lcout => \led_blink_inst.o_LED_43_16\,
            ltout => \led_blink_inst.o_LED_43_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_0_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__4991\,
            in1 => \N__5086\,
            in2 => \N__4690\,
            in3 => \N__5174\,
            lcout => \led_blink_inst.r_Count_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_1_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__5175\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5135\,
            lcout => \led_blink_inst.r_Count_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_16_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5036\,
            in1 => \N__5090\,
            in2 => \N__4994\,
            in3 => \N__4687\,
            lcout => \led_blink_inst.r_Count_4Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_12_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__5089\,
            in1 => \N__5035\,
            in2 => \N__4681\,
            in3 => \N__4983\,
            lcout => \led_blink_inst.r_Count_4Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNIGBEE1_23_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4672\,
            in1 => \N__4656\,
            in2 => \N__4645\,
            in3 => \N__4630\,
            lcout => OPEN,
            ltout => \led_blink_inst.o_LED_43_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNIH7VR4_2_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5200\,
            in1 => \N__4813\,
            in2 => \N__5266\,
            in3 => \N__5263\,
            lcout => \led_blink_inst.o_LED_43_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNIJCCE1_2_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5257\,
            in1 => \N__5245\,
            in2 => \N__5233\,
            in3 => \N__5214\,
            lcout => \led_blink_inst.o_LED_43_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNIVFIV_1_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5190\,
            in1 => \N__5176\,
            in2 => \N__5152\,
            in3 => \N__5137\,
            lcout => \led_blink_inst.o_LED_43_17\,
            ltout => \led_blink_inst.o_LED_43_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.o_LED_4_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__5109\,
            in1 => \N__5034\,
            in2 => \N__5113\,
            in3 => \N__4982\,
            lcout => \o_LED_4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_20_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5047\,
            in1 => \N__5079\,
            in2 => \N__4999\,
            in3 => \N__5098\,
            lcout => \led_blink_inst.r_Count_4Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4939\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_17_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__5078\,
            in1 => \N__5046\,
            in2 => \N__5008\,
            in3 => \N__4998\,
            lcout => \led_blink_inst.r_Count_4Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4939\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_blink_inst.r_Count_4_RNI488T1_12_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4869\,
            in1 => \N__4854\,
            in2 => \N__4840\,
            in3 => \N__4824\,
            lcout => \led_blink_inst.o_LED_43_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
